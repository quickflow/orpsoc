`include "timescale.v"

module vga_model (
	pclk,
	hsyncn,
	vsyncn,
	r,g,b
	);

input		pclk;
input 		hsyncn;
input 		vsyncn;
input [1:0]	r;
input [1:0]	g;
input [1:0]	b;


endmodule

��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_��J��≶���j������f����v��X��#Ο1�v�S[�T*]ZZ�'��b�&���\�uQ8)����/3{���>Bm0��̳>���T�d��#/��[r�I��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�PK��	�s�W���H�����_$
�_�{�=C_y�٬��$����?�\�+o�i����,h;��#m�����7��D��}LڳܡL���]^'�ie����aW>�m�f!�������IuL�X�������Ȁ�nW�4w'3׉0�G岴d)Q}��_>���/hv����!�[����Q�X��k��z�(ȗ�Q�����d(}����x�}'[SB[{��z��Sv���˾K�^= �J,�!�@]�+�J0:�yfJ/�a��V=�p���
Z�gvT)��}��8��p��w��)r�KQt��_��Ǝ�/���MX= 	��j�~G�-5�g̹���17J�_r�>��]�L�#��~^�&����meݻ�PT5����`�X���۶�"�m�ˋVX�g̉b�B��ΰ�O9��"uD*y�������`(L�)��w����;��ODK0���P�B��D��A*t��-���c������E������ŦNɚƑ��.�ʫ�^:o�]L�l���8��^�H.�zS�l��?#L���'�_zf3k�yW�� ^5,�9	��2��i����Fq�Z����W�����0�֖��^;���,[��?�h�lA� #XB�͛C��_>�b��L��}���*�A��m��=Q1}]��:)�=������:/�c�j�`.~F4ٍ0�������r��[���Ȃ9�?�I5��|~��'�M���WQ��l�'(U�(1�Z� M��g/�����l��H���|@�@�:6���J�X;�b-��raRj4�qH�9��U+�y7�'�!���p����x�a��ʄPzm4p������}�k�ۧ����0ߩ��� �ԛ��01�S���8����'�������������-|�'V�x��h`��,��(���ĝ��G)�e����c~7�)��oٞ0���5�B��Tmŭ��������V.�3�;#ޖ�>z6�]s�ӏ/lM�ӣ�%�KE"�i��<��M�~D��:����n�a�Os:���h�G�:wRW"$� N[��U��H�(g;;@�% �'VC~\b�mO�S3΅��o��x{.PA��f�ف>�i!p�lz��K>�ft�����#x���]�Y4jQj�ޤ���N��w��_$x���*���_Y����Ԯ/n��n)_�
���t�����$���(5/��_�6��gj���K�y=�F7hQ	PP��;����� ����>�"�WP�۶PD0\���g�����ѐ��͋t�P(�nU��N���r빋~ [��q}�SC�=jR��8<'���wNs#+�|�S8�L��Ѭ/�.Ձ/���A�S �a��@#j�?���F�D�Hbf����CHB��V�h��-~�&�K&�9�1C���6����v�V�J4���䔄�� ��</���������l���򒽨����	�"��!W���Ȝ]e ��T�s6;��T�ْ�^�^Kɖ�������7ؑ4�V���׆[t�:�IP�P�x� �Jy[�x�jdo���]�Wb��g%��(���H�(��˚��!�G��+�N��ԟ�L��w���#ê&
�a�_a�$;%��M-�rn��
ZG$���=���k�u�-�!H�?����Z���)g)�nV�eC�'�|^	v**8�&״+LΎ��0��`��~{��[C)�R$і6�
@�{�|�rO���H�r@�4O��J2����x̇
�cn@F=H�{ )�x���\�I�Lb� E��#V���2�tH��6��N�<���X:Df��ܜ�kާJx�����n�JCc�m�+ˠ�����\31\����`�=��ݐ�Tz�� ���]m�Lpvx����^�_��m{oh����3;Lc�YL���7�5�&g8M)��� �r���%�h����^_u^g�9�\;�%��� ƓW\}��1F :���'��:�����7���#/+�M��G��M���AW�E�[���
e��Z���uN�^2�d:�fsl a�Zm�I+`b����On��W%Qay+#?y�E�$S~�A�mPo�׽u��X1��?B&��OZA��44����M<g;U�f$9\Ĺ�`D���c�z*��0L.y��|��f������Q��w+At19��5c�̟��w�[�7u���^����W
=���I���� ��Ĕ�f��;i�h%���U�ړP^q���4���j#���܁N/i�؀n�����S(њ��	��D���`Z�fo�g�d�D��Q�I�������$ݘ+Dm�S��_M��ډ��J��Up(Ö�Dskw�$/ȏ�L0�~.T�\-CDA^�;V��#lF�$*�+��������M(���A�&�RIP���?��vH?��jj�=�=�XS�~�:$�c��ȑeC�C�����?
ݗ�u��:0{d��
��\-��?N���k8�y�0�ƌ+��N�W�T����n�ӄӷ���3�>���ksp��;�#�ڪ*�l���s��U~�1.�S�6+n^�d���6`=	$mT���Zj��E��a��!iW��N
\P�B��z�s�3�-J:��:��`JGX���=����S�M���8�)��%l�l���r�:2s7����Es�ݫL�L���86f3�b��:�7S��E@	7�ͱ�X�!�+��6k� �ܒ�d�^��y��{�iv���������
QS�[�=��ƚ�.�EY��?϶�ΑX��c ^�[zU��ۢ��2A����Cҳ$[�ԧ� [�4c�-��@|v���Ɣa>+�y#�RA��J�)�s�{|W���f��Fs���\�d�	��%����h9�"�>�ґ���'\�i�*�A�d���&�֝e}�.�q흜�85\�7se^�@j�W�_�)��y/k�u������><�j�izS\ABb $XT �4���/�kq}�wJ���K�R������+���P����Z���� �K�����K/��a*f3�c1r�O�D���-ւq9��4]���9�Wx�Tb�Z�q9R�JK-Y������u�w�=��Ѿ��b��y���g]�4�YwXEy�%�	��l}K%�8B{�>s��k�D_��e��(�����&���du[{^X�ZCăF��f�PMW����o&r����y�ԑ�2�������)mf�8��:/��ܼ��(�O��c�-Uv{o2�P�!�/�ӕ�=��&�8>�֟�w'BbQz4	cl ,A�Њ��I+�0H��M�@�[N�U����z�	��ژ8��^���<=����K�����fNl���p�h���,��R���l�yб�/�� �H ��<{�8X�̷`�K�{����o��mh�6jf�
;:I���1Q`����S�G�+���X��K�U�c�����\<���-��3ג�'�\��%���m"|�9mE��ކ���� d��؜F}���p���Y{E���/)w����}�c�a�H	rB��$���VZtX��V�,5�}��AN�w��:/��.n!@��{'-���v�6���=䋹?��G+t�S<��a��pC���I�e s�"䭱NJ�7����O0�ZPX����6��+��Ǎ8G:hߴ���mz�.E�� �ִH��j��)H�9ت�˄�YA���_V�m�i����6g��)��X��C ��ƕ���^pF�W����6��w���}�|��gm�e�9���dr�i�8&�*fA��si����0O��"�V�pi ��&g)�������ӝ�yruA�
|_�:�L��Y��pi�0~�ɔ�U:�|���ء���luͬ�줝�9��k���2��c�����Ĳ�zT��ǁ9O�ꖜ0�&�ߛ�ҙ��5����ے6r�Tl�K��@�*�d��I�%ǋs�7�4C��`�깐�V�5#�w�WN3�٤o8ig���(�5��fa<h�W���(m���a�ӼQr�|P�b�*�*�k	ugk��X���1�#Be��8��][ǂVn��w�?�ֶ��>��}}�ҥe<�m��+Ȗ�8�:
rَ{O��(
����"�) Hgu�*M�5��"�;2�`���sޘ8]�h�:�I����Z{t��*YX�J&O��+Q�g &� lt(�u�����]�(������G�7�/�ΐ�~0�Y�I�j�}ۇ�� ��L^V�� �� ��9 �}�:���_�����M��2P��R�Ml� �C1?���GS�᢭����D?��꜍_�p��$�s���;���N��WY�m�q�����cr�o:����<�23Id�"��RRK	��g%����ޭ4R
|��i�^^�m�%������ӥ��\Qc<	ox<0�� ��E�f��^����I���?B1�ƟNv�&i�-��"?�/�#���Z��z��pU���Ϩ1�r�(qL*ΐ��|���y����#"�����7��KL{c��ժ�ҮX-e��X��������
p	�����d���b�i�����_'mʫڜnoyG��jB���䭯�����,���uޞBEp(��Q���3>^EY5���}�2H[�+H2�>'b���R���ꪡά�n��āQ'���*�֑*�����~�Q3h� n\b��r�u�̱6k*��^��r���Ð0��7Ի�ͬG�K��E	�u��c�3��9�j��:��+L��|���`�
�kv5Ręz^��b��{�4.�<�XAAF`ld�%S����K�������4�3���Ps�N�>r�j}/JO�`�*�!]+�5��QҲ��I����܆��F*�Eo�� ��3��7��{��K����=���dq�����?��R��)��HS��E�g8��ף�{��^d�SU�U?&M���,}D�H������c���`[� �D�[2�V����ν{�����&e[`I¥W��(�e��9�˽ �S�=vڄ��x���g�Ʌ��{�_�����Õ�DM
��<1]�u}���-����+&�
H�Q����!�G=��`��q��Aͥ`�3X/Ŕ��m�_����s3��U�_�� �V?��N���ֿ��k��H^����[O�6"�}D�o��Y,|7
%��.�K;r&|)>~ơ$2?)7����S��_X Ⱦ����Q������q%�Z�)J<=���y~�!��k�1��E�1f����(�g��r��Ó�-��	p�N8
��[�'�~��(fȂE���) K$���?7)���ʪ��{>ԳV�ę�4+0.��땵P��%�E�Ӑ�DE�%j�`�&9M �m%��?H��!
1�7*��ؘ���L��!wq�m�6ʁD�}K�l����,	�����݄tXԦ�M��[�;��}���ۊ/���Qd^�h�����bA�ᰧ>�/(�)��2ň���#�����e�<���r�w�����kHnß�ԟ�'xv�4nw~�	^�1ܝ�4��~_ېp��C�N���YPs�ݽ���D�@*����UkY=�MM���q�(��ӕ�Yh���Q��P�o-���E���m���<C�o�NO��+s#�kC�l���<\�>��.D��^e���ys��b#4�Ya��Ugͪ5�_rS3��r��1�e�@�	ԍU��G��|��a�-�: Q�ߟ�����2j������s�cA��/V�t+���3-^�&'��:b��ϯI�m��{t��������ڰ��Im1��k^E���]��&~��g�����Vg��ld�z�+���l;����ťڷ�{��_lr�t�K�v��ӱ���Z�<�y*"8:G����*����٦YG���^1�՟�H����B��A�&T�N�b��7I����i��T��m�j)���0��i�?U_�`hs�Je�l�΃Y%C�9_�n"��[�]�cI����4 �ţN�0�����A�&�e��CS�0:b���lo�B��uZ��Hȣ�)3���	������ĪV ��Mk�O��Uڋ��gW�M�M�(h_���=��bn��y��'ߥ�"�vG��!�*����Ж�.�Ĭf���D~��"!�qO\�$���/:W�P��)�	�˗S��aCJͦ���B�h E�� ������&k0��uk!M�f��r�d>�t�)���N8IUl����X��>��'�y��R��a�h��IR'�#]苏�����&����S~ZkL]�V��h������NS��i1��"t��Ij4 #�K7����s����ւ��T0��&���Ԝ�Jh�����,۠����J�`-C�aゴZ��I&#�1��=W�c����e��5ć�>53���J���F.r�j���#�I��ոg��vf"9�.�-�{����s��1����#��X���A���Di�fK�[�
������3�N�$d{Z�Glr}�U��S�3-_q0 �|����L�*�����ߟ� ����C�N�6J�����
(ko����Q�&,J[���oAb7ڕ����W-f�$Y��[�F}z���'1��_#oRH'|�=�bx��@���^�U�v����hYj2�!��wf-7����?�b�M��h&B<�aY���ά��t��c�^�H��Bn��>K�O	Pk�D�o!)$�p��`�����h����ˬO9郈�?�{��+|{���C�H��3$��8x`�j��x�b{C��t��5	z���y����@Kċ�)�1�}�5�DU���Z��p9�k�U�&�ƜՎ����)�ҧ�����Uo�ӹ+tח{E7���A�B+4'e��H����'���#e���5d�ZP��WS��,���9!�/��L��wP�7]�{�N��%)�����-����`7%xO��7��1y��M�+�M�3š��D����:�<�esoFq��NM;�7C�߮�~.)b�A���?o?#�"t�;}��>�Rգ�ᔃ|Ǿ���`,��9�Y3o��1
�t23��Ć�q6�)Gɹ��ڦ`xhR�KK�=۹�+c�3���Sv�Af�&�][���13o�u�Դz߿�֬.�0Nh��w�r��M���V,(LV�q.�le-��V���S��Z�bo7e�7�
�q��2���窎e��屬�/������M��n?���mU(�^��#.3D�j�F��t�@#��o+O��m���_��?}���.ۉ��`4_g}�A�$�	?0mʻ8�M�Cz������F2��W9R����Ƹ�߲Fv�$e�e\cB<{�����<���/YT����o3$'�����<����E$\���[�h��Iv�mF�W�RM��K�J'��H��	İ�#+�{4���l�hx)����|�| >P?M���������� �ɧ-�l�wh�!�H}�l��~�K�♭��o[X��A��A)b��즵�Pu�M�8N�Uε���mx��o�%"�w	�<鿇�+
��8���ݐ~�W3٧Lm�d���f ��>���;'=[5�����է�ZFة:�w��m20�A�a؇y��\�� h �u���..��`}��F${p��Ͽ��x�
��:dvC��S���;%��S[G��=�a&��NW����V� �x��������q�)+����n�凟����؉��s��ɇS�׫l�|����!&DKO\a��t�����"݇s/���x���j�'���h��w~|�y�h���,L<�'�%��H��nx;���j�.�O��^?�Y��`Pz�¿�/���Y��E�X�a�
����C����H�mEg\A��pBv����(�6���b���i�0�@�j��X5O@�w�Q�ɛ^��
_��9ז��9��8�qƏ#j�A��vW:�j4%zs-�Cbڍ��7{B
�C����
^�4a��é�`�=�ʎd��.a�e䖣�&?��r¤ѓ��t���)���d�eKlf:�з�y�lM,`�A/lsD<�e��F�?���ԧū����D�Z ��x�I�	ϸ�nl�
C��N�=�,�}zv䬡_�r⪃TfxN����	y�P�g��KU�M�bx��c���!l�ه��_���]��#z���"�C���WO|H1q���@*��$��y5��K�+�u�"��RFB0��"�$D�M�x�磪�R�-��A2 ����,�!��F�fA_K����/ǣ�>|���#`7�������mǚ�z>QN����_��/�q�%jo�� �%��=��fr���^n��v0��ej�v���p�/ע��19��N��5�SD]ҙ��|l��g���&=��`���q�YM7~2���
G-X�Im�myR;�l��3��K����{]�L�+�Bg񘢢T��Bo�d�`,�Ne'����!��f�C��֑�Mf&��ǈĒ�T;9L!�h-���8�x6�#�}1z$��Q?���6�"�.U�͗t��~Nh��&��P�"��P��3Hhjk+����}/Z_0��/,�B�˻~n���C�K2>�ŉ�j�.�aB��Y:�[�_ͯ�2����N�fn��2��q�*gW´�!6��Ae-������Dr+�I]��˾
��`&��S]<{� {P�/�)1P�Hk%�6���Qq�<5�r;��./�Y�	�>���lG�����J��13�\y� יh�$W9tSR�D)�צD<�Y���``ir��,c�VW�4<:��rեlO��������aD�HB9=	N��2�d�Ѫm�j!����P,:�C��W�6����?�D�:!4Q����U��9z|p�Աe��X�1,�V񠙒_�.�D��5���.��Ac�4�1�5����(�d������Ul�f��f�K=��]��تi���HY�Gz;�B�wc(W���"D�������C�w��n� �QG�⦉��j�!7$�}�Aסg�U2����m�.J�ܽ�;.��#��Ǝ���_ŵnݾA�����;���z��`G-N��"��_���Y��l��ȯe������g@�s�mI�'�ǧN����y7���r䒵�p��n6Qa��LI��Z:��W�����TU,H�NS'L�z�<z�]��lS��T�ܩ+�����K����b�7����9��o6�\Q�a����	�8�LӋ��X�[ Hai�7�{��%t�ޢ���	ʌtX�݇��p��r��V�-���N~���'ݫ��U��mB<�1��l
$��D�\�c�į�)�'��L���+"^�|�������nX�b,w�j���o�q���)�G�mp�6���ے���y�娟���j9v��N�	��׾��,/�� M9&��Jq��!1'�Iht!���wCP���A]�v���j��,U���|A�H��e\�6�~�F�Ƽg'����+�k���]Ch�3�aj߿��<������6�5��CG� ��IF�y�~�L��٬7�}%�F�Lq=�D������Otk��2u/Z�@�#D:�~�O��4� (�abW���k�T����0�c@�Y�]���"��@�i�g�0+���>��U����]y� ��e0ߨ���"�Eز��?dG)9d�۞�Ə3g
������]JX��:���R��ZM� oG�K3\�YkvM���a$�UԒR�?�o#�����\O�w�!�j�ٛ.��T��+��^�j��^��ߏ��}��*i�1Le������Iu@���@� Ь�����?�$m*��X�*q�V"JR=���a��}r<w*�I�dN�-[��5	�<�tT����X��'ɑ��'C%��RJ��r�C��ZQX�=w1e \⩐��W��Y��	_ؚ�Х�a�l�rf��(�S m���y��q��B��ΰ�7��nD;<-���2SE>�l�15��e}�v/���V��b�[��ۈ#+�N<��}�l�a7c�)� �'��X�i�9d��������� �;=|8�E�ﰞ<��0� v_|���ȇ��'�c����fL@����G�	<�s�Mm�w�K﹝�6
A����kܥ��&�:�D�:N �Q����~<�Yb�\o��Ui��""����P�B{�&&�i\59�c�F�`�gV�$�M��:�iKLNкX��Y��^d��ɡ�(�o�_�6�iZ�}������q��~�o�tS�$�/�� X3���0\�~\Dq.*U۹�� ���%��E�k�M�5�m���MU��ү������H�p�7]���c���z��}��o`B�E���j4�ƕ���� �?����O�!a{Bf#G	���K������G!e����r�W���\y���=�"}-���r`�GM�*,#��r��*����x��c��������!��3�.[�x��58JMZ$Sa��}��<�>�����?A��S�r�V�0��:��d/��.q��)0	��E#�2Ⱦ�s�%�fH��p,��N�p*>(
���>���*���o�3sJm�ml�:�� �~��E�*�R�cf�-0����Bir���7d��a�Q����MW�x�NT)�� 1qRz(;Jτ��P�hѢF"����*đ�|g� 8�;�k/H_��-�ߙ� ���QI�R|m_[Ȫ��ɱ����H�X�2'��"�Ɯ^��b�� WrS�?�Bk�ݲ��%Ɣj�%�����J2J/�6
��X���ň�����������-PWi��cq�bJK�\�T��i.1π)��P�D'��xaOv��$�7�������t/ŝ2��x4�κ�d_�_{ztک�D0$K'{b�zgPlx�����j�=����Gh;6%�Q����G��u�}(i�� ��(W��l���ڧ����iA��)������j=��]y�⦅�S�q{�~���Q�������Z�u�C�2�Sӵ0�L%mh��A�p��d�� �	�,,ƒ$�E.��:�� �(��j��� =;8�i)�H��.2
��<��AHmh��ʗ������]�el
�'1�&��oZ�vvT�*\���
񆠓�b	���m8	��W�k�B���'hMp��xuR�f^�����G����нC�΢z�2�����r��v��h`z�uO�P"Wh%c�`
����2�0���i�O	k���+ф/^L�=�#yk�B�Q�2��|9^d��� �=��t�h�����T��b��V�[��x���f�>�%c�St�7p#��5*ƋF����`�*ɜ� �/���eA��_��&�k���Ns8�a�W�ǳ�d�D-�2B�WM%�kǢ�F+�P�u�������Q)U7�-g�lX�=<����zc|��Bd�Ơ�nHz�B��#�/�~�3?kw��©����X�c�[5�5�p�f:x�IY��s�My��c=O�����GX��5,��#9�QՂ7f��/,���3���ÊX���k2�x����\� �B�����b� ��G�B�����ʎ�vqC
-���)*��|7�M����ch�xD���j�)?��?�I�C���:*аG���w�:S%��d�\볁�p����/ة�[X�Ll��2�El�F�2)�	]DB�H��`��~Ҏ#��L3V52�pH�n[���{��U����\[���}��~�[s�{���^�DV�a�����t�W
p;�%��0�&�"�d���9fv����2��cڵY[�gn�ύ(��.�H���JK*���y]���0��Ceyp��Be�(��EвW*'����c(S�X��-���O��QG�P����������~>Q��XH%�͈���ع�P��]ƆMt��n>((��}���s|�����`��[�!%.6�����7��g5B�тM1�+�.����v���"�kʅe�ȝ�p.�>3|�+�DΆ`��'��<7Ɠ���=�G��G�fuTƼm�I����C��,�P���5���1Ǖ�_���{p�reZe���zIQ��9N�[#�nKbq�R�}������~Y�̆40�Q�f��l��g�A�U=�=�FO��;~�,v�e:��p�dF1�RI��R�(�^T�(I�@Q>H5s,a�xX�j�
#A5n���Eʹ��j�XSs��JJ����*���:��&4��5ye�si�ƶ>�4k��wè�ȩ���#�OM|���>�w�_�=��	Hs���_�@$*�ċ�heq6d����xԚ�z���㾚�N���	�'
ט���<a׍-���oyMOjf���S ��`�߻�|��.���C���ӌ��rB�8�*�h����Ƙ�o����N�ԅz�dU<�[�/��nh=])���%�a���)%͇��Y��H�	ڜ�ଌ[�c����0\?sb�̨(�PM���)���jZ�W�%���V} ��sU����Ə=]�F���� �����=)���[`G-dS���E�'&������E�K]Ƹ�t�0�+��ʵ%Y���!gja�jD޻ʡ-��6p�Wl"�w�6r�����r�?�_�6�l)�_�$�J�藰��yUC_��S��t��X�T���SY��
��I�(�e�It����\h�l�l�np3Yڭ���J�͑���Z4���l�L3ʣ����	J� iα�`�JqK��3��d	h��
�=9��f	��Jj�9�Z��+���f-��-b�Y�)Nf�/X�+�x���&���z���p��қ�)��������\�jz�@�%����tZjھ�ۡ}1<�tu��y��ԞW+~�Xmh�A�>�T�f�{��^�� ې�тI��Ԃ��J'�&<L����ڍ��U��R�����0ҧ��#��-��ab��d��|Σ�\��r�3��'M�>�jmK����Wk^��H6��C]l�)ì�{�/�X�K���������J˧�;� +���ӻc�.�t�G�+�1�*����1;L��M��fM�����&�0�L�ьb��Y�t8Z�(����.��B�TwIPJ�0�rܕt�X�\�C��t�o3�=#������ލ ��]��������@�<	�v�ƨH��i��O�p|�i���������Qۮ"�1|�*�L8��|����½Tq�rf{����Hј�c_�ױ�x�QT5h{�ps%��3@��v"�����;SuH~y��l���浠�]��A��X�q���Ͽ�pM�?��8��?���a���𠉺p�{9�3B��^�q�� ���ы�Xl�8�$�Y� ӣp�(7��ı�s{c�ʹ�r�N)�J�\�xB��X�����if@�w���|�?��8�󔭝�Vx���y�\��Hkk���n��o��,���z$|����ɀS�A����*�.��d�*8A��s�Z`� �����E����?�A^���u9��3������y���/z��$�����K��f����=Yb&	y���]A�����EЖc�D�-m�,I,��,�$HI�G�.<�N����٥?�mh#qre��JUP
0[�Q�5|����	�����n/di��xW�����*��,�H1cn;m��sAq˾t�9��#.K=�p#W)��a��o�r��f]���/���w��#�Oi(�PX�H p)�؍����>�VC ����X�vN�ѭ6��'T�Lh졨�/0^���I�/2�}D��!��I������J^���2Ԯ�CZ��Jܒ^�!N2OBH`:_	%`肈�C`0�g��D��x�LO%j׆��wy��F��+�<�&�Q����Rt5g�.iLN�,��^������B�d��r�Za�)�`���ҿ,��Y�`�䀠>���꧗2�I��{g���Ƣ��\�������y#*E	23:��@u��
�-�{w��[	�γ�o�5��Đ}X��T<J»E��I�ߨ
�g���]�AHA
?�Z���/ӓO��H]h��g�:��w�U�f>���Zp�c�s*ė��:aA�α �A2�k㰸�e|�ͦ\k��k�k��.��.&�Ŷ����o��vQ|76��Xn�j��ߏ��$��p�ϡ�Β.��֮'���$j���*TC���,�OW�NT� U�Y�ܲW�:�x�_ֽF���+@��9,֍+dىLa��q���[XITg�	�!0^�2��-|�P�#$2����5uO݇���N�Q'A����*���z-;i�q���)���P� 2bO;!���f�-&���˱JT���9��c�O�AL����;'#�����⁣�p�b�wA��.��<K�!�7G�`�蝒�МVA�v�� #K;@]�މẆ!���ȯ�?!���9�϶��;��E����/m[\��]��iـy��ze=3?%��턲f���%^��20�8�0���&YM�*��������Y���J��&�&�Ay@�O�;8TRz��y7�d��f�� -3D��uO�}�G>*�g�Zg҃�l��u�|z�ڱ3���N��K��3N`2����=���@o�Ѕ�;��:2�Cf�5���>~���u^=Z��a�������|��Ŏ���{8@D[ �sw�㊹�g�(M<�.px>�K-����h��9���BkSp��R�\���A=r��{��T����3QL�3�^��NA�*K�2�o%��X�*�����F:+�V� ۨ@�v2����*��וe��Q{�x,Q��p�i�z�ڈ*f.�|K&Uk�AY;

E2�ԋ�[��B�=�%�`�Ҧ�sو����i��ggw�Hv����C��BD��#�z���w���xlg�c��W{��S@�[��r��Y$X3{��V5e�;��az���7���X�&/I�5�3��E��.������nX�e10$5�=$��k�$�l���rG��&�e
2��߉�0&�Q����yy��"�4<�L���z��U�K�?O9zn��H#pi�����b/X͑�]kn�`�f���BH�o<ru���M[�;B�輩�չ%v�a׏�E�j(x'�M�� ��i���R��Ut�э~p�?�
������pi(��L��ˀ+ޯ�y�d)^�=���v�Ŧf��12�e'+R��x���v]n�rl�7�k��2vjy���9$o�2���7S��ّb�z��n�>�Y���s-�6��}�c&��cF�זAݹ�CBs��d}唇�=����/곟�d��H1B�l��L\�s##���b�۳�'��eFbU/g(�����2��Wp0����P�P��O�^_�sC�){�w1'�m�&]E��s�-���~�y�b���{MZ���buE
c�zT0~w�E�n���E��(�U]�J*�s�H��J2ķ��{־L��7�t�ce�@P>���/���L
��n�QLs-B��̺��^�Eqp8�J�Ծ�og�5;$541��i���V��f(lRlP�%��n��1�_��4��z�"�S����P��jl��޳{2�?B	sVw~+�J��H�a�#�<�ם�Q��!�7��a�X5ir�j�L����U�(��9�J�5U�]����BͧG�����Yd1��@Evw���Vnl�|�Z����9���W��;$i�ցh"T�6(�?V�9;툯a�����QO���/�m��oY�8.��Tf�$U>*�	J7*������kw~�e�f���G�#�;?䧋�[P���P����p/�)g�4Uxp�=dO<���o�f��c�u��L'#����}��N�3��ؙ�я}Z���`������`Fp_̝�2�
�o��ш$��R�����&�K�]�mdo"�� ,w�Z�\g>�/�3�"���<�yϯP���x�d�0CP�)X�z'�7����Eׅ*��-�q��n^D�����&5���/)�j��F���e�@�1���,DF&�틨�ؖځ�i9��?��(�1�0x��O��e�!CeiJOC�8�,���m����p����J�����em�.���/�=��M�n��4���\ou�֢#����W�;��b�Ԉ����wO.(Yd�ڴ��} �I�}t�ub�9��
�f�(��L����O���Z��vo��l:��ژ��%@�b�����5c+��&Jo�+�*�KI�*��:a�FF�$ǅ��0��熭8�E�+U���<"1�e�3�P��g|�S��i
+q���Gǁ��µ4)Lv���W���5�ks)�6L����TG��ʥ�� �qg�;v=/�� �D��;I��ry�[��������!r:����v����2uo A�k��5b�?'Γ�#9��p�QU���ڌȮb��v*!��1�9��bºMt�u�qht����A'��'���1���;'Q�zT0�X[3[�`��{�/nw�Ű���Qe�d��Zy�v�*
e�i_�EF|� ��S%B�;n'���ysQn�	� +x&�8P\���IS�����X� CI\�KZ�(��4 �`K�8�M��S�l�G�\��C��B�M�W�wv
�6��f F�]"0����M�u(�q�^�Q�j������쏚��b�%?U�c��o�֝�UE_e���},:�(��O�L'��[G��"�J]�J���U�T�4�5~0��z�6ܻ���K�ͧM�2�Ƥ��ά~ִ@�UA^�n�p�S��Cf�d��H1���,�V��y�St�9�C�c�v7!ɹը�4~ �������oU�7�1���u3<��/�J� cNa�r��I
d�XL�\���D�/��c�ޡMp;4��`�{4`��B��|.T��Pz&z7�K\%;`3|�+;�����בk'8+�2�s�����>iÀ��΅��C��^b��=�` &�рRX�3Q�l\�S�����Q�U*��"��w{Z������ޟ"��-f�~�4q_gZ�3��1�����3����\/�8s��R(��	���(Ɛh�QZ��GO���Я+�@����^�=\��n�����Xd�ϴw/��^���d��^h��$��&�Sz!X�1��u�y����b�v�/�|R�2�ww��f}�uqɜ2�-b���P�	�f��D*����Yip�p���S<�b�XP���(T��_]
A؋�ϧ�����\�,�0��8���"_��y4C}Y��Tr�C8r����#>��P��q�薼�� ��1�����X���GuI���;Q���$R;��)�S%�ϴ`=�KNA'�|�0�L�l�6ir��������l�X/�,*n?�)}�GO�D�>.���R��a��>�=@�yJ�K2��H��+9*.B��x�Nvu=GI�Ȣ������/n����+�`t�Ǒ�o������9�ďؠnh��M�!��m��y\w�¼�M=_��JOH��<�C7�Iu��h��͈K!TF�į����.�|����^��3�q��D�h9�~�E�gF����W�XӐ:G����"�����^��(��C�^��%-V���-��ҷ�f��d��do��pK4�q���[��y�$Tx��qpK/����зU�^K{�MAݓxr�����.Җb�}��aZ�C�Z����2����.n�.&�R2s*%J�P�݊�&������x�|�D��'�Pbq��LH�+¸�7�����!a��0`�_��&�J��+��GFۯ�5��(0Nc�U��}!-1H�����'�xZ��Q��R���>}s'����w8-�Q�g��e���9��hOܝA[v�oJ ű����Ti���V?оYJ��xrS���1A�F42=����}	޼v���N�r���D|�>�j��T�k�%�N�Fg'?��v'\����ͦ"h5(�^�1���)��˄�d��L���0�@}�gI�%����r�J�w�j�g_�ǺH�Z�B�K����ڮ�8$R~ޞB@��T��)��'�-��}Fm�|���tI��>цX��^�nW��C0���0V�}9^X�6�aLF}�e�gd $5�4aZ8�T�0��{l��_�{����Qꍤ�8�=�n�0���	��0�x�ДV���V�2��{z6�2А��ߔ"Ry!q����Y�R��s.T6��0�x+�ԀŻ��K��j�*-H�%J^o��_ƉN=�*���$'�G�l~k��O���7��UY���]wze�y��*���X�6��t���$����1�k����Rx��p��;��a��fen����^�Y��˒[�<p��l�綊N�����^#�C���x}�����;�'HPlt� L�{4=9'�XG2b�+���<��j��v��B��m@�Jْ��"�L�}<C'�9��L����嫷p�0k��"5/{��A�-G���g�V�V~�ݰa�c�ja��E�����9: ��p��sYs���'GQ�/��~���j%S�Bqͯ �m����b�&g���6fW� �ob��%q����c\UE������P?ɡ4�S;���<�����>$|(��2˝�\l_t������q��D�z�û��i�i�`h:D �fQ O	^�A�`Q���V�_ўJrW�*��q`څ:�NS��@X�� ������|د|J��_��^𫮀v(���Nq����{�q<%Mb��	��U���ш]C�q�{h� r�QR��F�
�pxa�y��'BT�����[����j=��,_�)��"{�h��8�Kkox���5y`��C���g�Ԓ��v���0��][m�fCu�QQj��`�!;(�Α�`�n4�����b�%���>Ӻ�2+W�D*a1�L�K���ϼ���r:�O�~���r#�CEC���������-��ta%��\ح�&����8-Y�/l�s��h�=�3�a�+O�Jα��6�~��H��v��Ȗ�hXkLE���B�|�����������_��u0��L�㻝���D�Hxk��x�_6�w����%��'}7���7G��!����В�� ��o�_1�t1���q��#�&����
�(��)����FBo	
����*	������ex@sD��C����õ��f6��ކ�����i����]���O ��L'�-Ė�,�Qww� T��692�u��
{A�����%��v�W0����":�߹�Ӆ�탬���1T��K����E>�����M�)��M�L�}�:��63[L�_����Z������ܡ��������_�H�m2M�d=����M�������1ZVJ�(�4jhPz�d8Ɵ��@�`���D�b1P�&MG�txED�r�;��#�>�q��]���~�JU#�D���<t��e�cE�N芺����w�[�K>~�(W�.]@h+�p��_�{0��P����0s���5�RW�uD���j�2N-�� �-�s�GW
'����	����O�/�d��4��YN�IC�S0>STRks"��ˣ0�FG{?���y,ӱ�R>�K�]���ݠsV��ʊ��@tY�ȼ�劯3��OhE��&zn��EwA5��.�8���x�Y����l�_�a�<�_��EFLLѳl@����J��XM��5lU���-͔��P�3ԜmQ��s�`��go�(����]���j�V��wz��N���KI��<�����t�`��I �[a���j�����,v��f�yt?�-�8���+����%?3`��F�e@�Y2�.i�g3ah�ѯR����䛧����jp^���H��ZwΏkܛ���w�
Nẍf0s~fw��0��9�;����4|2�Y��c�K=W�jl�f'ZY����W��K���'z�G�~�)>����T����F4��U�'�'��?>A�y��d��7P�>��M��8���X3�F�a�D6!��;��ږ����T?/qj�̫����I֟�u�������<�F���Ң�0�l(�c4t��*˓�L�H�<y��!t_��=����tc���[�b����ٙح8�������|�j"K|=�K,0u��տ�,TX-��)J����$�e�8�� �j���#��_��t[1}�
�T}�)�+�c��Ɯ��}q���Ђ�#���
�j�1]�SUǆ�-YK��>���xh7�ZMO��ǵ��c�ɐ9�����k�9��"�x����� }��.7�]y"?�aZTH���n<�T/��p42���%<��:M��?	����٠4�br7ۻ���0kpѥ��c�O񢺓3����k[�"�ϓ��ѥe�?�X��z�N��.�JzϷ��o�	m�*��>]�i�=_�@�p��؅n�&�$'G���{͗�0��҆�X��k�fÂ;T�`�p�c�4U��{7�/��5��E��f4�2�N��$�:{�+
�H�
T}>�⍶V^;WA3%�)��k�/�E�ҋD7�X)�=���a�-��Oƫ�26u/}��Ƞ܍oh�kG�)/C�(|����k'\*(k�v�e~ ��u���Ӛ��ޮU��Yd��;�p� �̉�Ym<�t.�}X�qѾJ�A���u�6���ſ�نP�w��Z�jS���� ?;Rq�o{�_Z<9@��qAR!s}f&�O�P:ͫz�Q+)�]�ABig�;�o2�f���M:�:�
S�E:SP�I�饠���@"�R��sG4�0�V���Z����7;�r�V,[{��w��N��ƈN$��Dˬr�D�m��e�����(:t�FO�5�V�NA��,��Q�Hn�#�/���,�������U�=���a�5�xy�N�c�Xi�u�~�5�_)=\|f
x��y%�������o�a��K��M�)?L��f7yR�h�����c���+u����V���ӪX�BOrt�n䳚�5�Z��§���רoA���9�}�Mr��~_���|բ"�J��w�S��4��/T�Y�Kf�|/~��l:���ȔT��MA݌��
|�ԕ�ɡ!�1@��*�66��-B)!>����tq�hΧ���:R�h�'��n�G]Ƅ��C:I�Ά���Y[��$�72�ӽZ������n��Wjs���&���L�e߮_m�N">[!���:�T����&s�����������9�}�7=h���x�����q#�gU�ZG!����� ���n�+�*\�81W�/�[ͦ8^�7�Y�
�%�����ȥT���A!���>!���=���D@�����T\nȳ(OtNF
{�j��KOV�U�(�R��5��zcܲ��S����!P��2ml�و�j�EW�?��5�7�����O�nxIK�^�i�w���JQ=�Z��F��!�2�i鰟Ss��#�� ,�);0��e��}��&�g�2��3���Vm����c\�9�����v�>"#��z(r0��32�zY?{��M��42G���C�%8�ܢV��sd�U��c%�8�j����eĂa�S�0�S����������.������!�B�TYd�_Λ��%�^�Z��\`�_��R�%��N߰���s���6��觝R�h����rF�������"���8	8&�v�9�o��6W�a��\[U�=�����.(�C]y���N�õ3�&���9�Wmo8�E/���@jh�	!�Oޗs�0q��/�h�E�Y |y������ ���e8�P`�6������y���j�]:����ƁW�N�D_g���m��Ơ�Ұf����o���-�����=�i����lK|�k���HFP6��ԏ� e�A8P�hs\�G~�M�2~]����Lc0�mB}���?A�ޜe7��Q�0j$s�$��}�}4�����X��`M�q3��x��~�E�J�P}�UV�%�ܳ���}(�&Z	�¡
��KU%��+�X"j&Lԉ	��͉��T���/����'اӥ���	�����Q���^����v簻��&0M�,<z�������Sg�ꟐI 5͛�� E/Nl�/֠�G +h�ҳ�������D�����W���<�)ֆD�#g���n�o[�:�`?����!:����iQ�숭���Ek� >[�4(��́7x��M���}��� L}S���ΰ���'�H)F��4߼$_ޟ��� �������#e�L�]�� ���7j�tK9p`�9j��,��q�y'�27�A�&��E�/���u"]��{�W��Fp�vO�⛁��!9������'_������J0'�F����Qt��X,` _�E�6�mr讎0`�=mX<�����R�1U!<0]��`J_���D�ΡFFs�aaw����\��������Ek67W~��}FA���x$e�M|�?v�W���2���X[ ��V�����˼�[4:�╊#s�]�?p��c%H$��;Yw\���wooDL��<�q�C��<��Õ��\��f:Y����`1���o�ِq���_V�#��\�	��VJt��ck_ѝKd)����דo��Xql��p&�8���n2�B����5�8�;�?���S5����S������й���丷�i�ʖ�v��I��ބa<�X�W�l�����(��dW�N�yp�N��ZK������-Qs4WtĤ�rpLA�W'!V��݉|4�n��j0�x�PQ�l�×�腪4V�J:�7`?',-�����8�cE^@ͭ��*f2�u��*Q}}B��I��ݤb��<�06��m��ߵm�XS�38v@�7�|�^�鈀찼�q,4��kG�%L?��&V��Q�/&�ǔ+|2�i�&"��Yb����A��6�������Q�@vi4������P�-���g]�A.�]+�P���PUٸv��M������*PF�n~��=^��᥍�4Q�S�G��ޝ�1���1�7q�rXu���o�E�K�61�zo��;���6#X��h��WW.	������S`"�܄G�e��)�2"J
uQT+*ܑ��u�ў���i� ��ֈ|�9��K�3H��g�_��<}k�h��(9�ԗ�8���?F�%p4h5�a�
����%o��߼Li=�C!u��׆�� 0x�7P!�M� 	M{�����7�flM��΄ⶱ�� )c��v��5�hl�q|*H�-��H��Q(�|{ԓ��k�
�`�̯�t��z@G��5�:�j�ov�+^�=�+8�(2� �Cr���}�?�y3�!R�&쳖\�]I]�y�g��q;̸�9k�2�?�����x���tտ/��|l^��A;�$-9�;�i'�w6G�`�g"����[L���x�������3.�%�Z�����^Sd[6�)a{a��z�������x�i��S!��W��&m�(�K�z��{l<&5 =�s�+*?�έU�i����J�lQ�ݑ
��ΒGH�f�����{ջh#�6\{/���H��o�E�H����&��q���m$�6�6�٠s�z�Hu�ϊ��/��1�4������>Cˡ>��S��@�vxkl�om�gA�0����
v����yQ��|�&�]-+z
�9֝6
�u��n�2m׽~ļ�YB���?��N��ö���ID�wd�����O�D��<�&k�)��F�k�үR�M��u�bd��Kb���<�M�x����3�k$BkOgl\�}$��_���g��6y3_sw<��"o���u4�%:�G�WsvW9�*z=�WL	�q���������ߔ�>�!Z��{sWP�䳪���t�ch�"�������%,��l8$���������rY��#O!	�}q��!#�߳]T|X�G6)���*�1t��[��9�8���
KA���#�x �\2����i�%һS��8�� =�A��K���/����y:�m$#�ཷl"�����2��sk�SMpG!��ч�~C��G���n$������e�`y� ���6Ÿbo{�G�_�`��;�XT���k���I	�9�G��e�ģr[1���0Ĳ��`��:�ȟ6^�DJ~����s�M4�1��-8.����4?@�sқ����2�}u���H������>�y�ٗ�=ݛ�6ɣ��K��2>;���v	�:}L�)X��h�vt|J�������Z�.NZJ2/��B�+a��e�	�hYD7�Q� ��[��ٵ[�h���V�iI��A��M���r��質%o�:����J4��K(vA��rz_ded������?�Wm�1��.��ze"�B��ғ�����K�揁W[ɟ<��u��|Q��A�_��q�|��\W�}~@=~��FS�C�����Fԍ�j��1.w.}c�J�3%�$�V� u��3��̷�bz�Muj��|)���D̓^k�gn	�n�P=K�M+�a�Ż��AC���T]��.�P
������"W��������&��0uH�����ٙ�~cȴ���o�)�4������ZC<�X�"�L#�z����i2d?���a,7jX)v��i�GFJY��Zj�OO��;})�}�`JC�<V�G��ۦ��c���.,��d޻qio�?�_N�����sE�_��	�L�J1J}��r�J^}�����ss��Ǿ�]x� �s�z���a蘘1F&�+v聐�$�,�<����OE�M�XL�x6��������N��g�_xC�m?)��M��*M��DeGI.�VwY�h��:m4���}��[^1���"U����`3��ӎ�$�ƫjq�� _z����� �Y��DW�`f�'bx�c�G�����>�*x0�<�_���=���{ڞ\q��:�I�+��w�9��Rh��%,lְ�fB�o#�DNhM�?�y��w�1�*,e|�8)S�'Cj��>�P���!��yR��Q<5�!�!�~mR���C:�\��ćAhh	�^?+�d�4��xW5�Ʊ�p��@����͢VGi��h�\�1I��(���3��P���/�膍�k�ޥ�ɓ`_�*	]-3a������*ȉ=u�����%�9�XP�s=���vN��k�"�������%�
��G�y�q�G'K�_�T�]���#�����	�n(Q��j�w(7�p4�ם��1G"%mx��^��Uyw�F��E�QH%������:fE��#&�Ц�q;Q�'R��d�˹V�̀�o^�K@��t@&�G7_���;%E�j�#s�����̆y�)�H��}�a�e�;��M�Uf���x/�7�&`���ה����z�<��s��@b}*`��ק�����o�_kE�*/{�/��ݾ�@�֤�t�$m	󊜉�U�*�$b��F�A�t�ˋUaK;B����y��@������Y����w,����ZV�e�5�7p�L��1^)�������P�܎}X�4����K{�1��Z*���Mk�'A����_za���RP�O��~�J*����i�c�k��e!�d_����k��u����lw�����k�R���s�5u��ZR���9ގk��f���b�9b���?X��n�7~z%��ݞ9{��
Lmw/*�<�CY-�f*^��������Ej��0WW��9&0�7-����R�ʀFr���瀄��]�
~���1�GΧ۩�d0H��}���sؗ#.@X9�V�xy�X	<��n;��Om���f!	O�-xI�J�;ZK-n;ФP�^�,X/ߧ��檈�?F��mY�8�بt;�}ٙ�NY������;8Cb&Q)��g�#����b��!�|?İc�N�*��/��t\��{C۩L̇�����YY��9"�4�ʮ$Jj�,�\�-a�_�˔����>��Q^�52#����e�j���o��cM��3�����o9x��]���'`OAe���W=�.��5m1��=��kr���g���t��u�S4UM��T+̐Nm*��yD#� ��������:C��Rv�^P��Z1������$˅��
�7:�=�^�&v�I��E+[��6�i�c���k��9����n�17@��!-���%���&b���硜4�%�<k�t�N�]S_��� ���i˪W���F�s/E�O�J�.���aU!@�B�p8�Kn�P�����ث_|�MB�R��OJⲥ6t�{�r13����Ǯ)�18��*��suH��T�@F���^�f�[���,�k59/�R����*���_��,O�x��E\|�8���`+���!�d��{����)�i�tâй�0}�c�5�l��ꪉq��26`��6f<���U�?a����`*�]JO|ǂ�|����{Kx�A�U��M_���	���(���~!9(՟Y��J�Z�6�|�ֳ� 8�ܖ]#�yM�B�&|�el�YUͷQ���s�b0�~�œ]��u6p��K��<˿Z9o��}�I�⽁�:��!����\�ݫѕ��3����	ѩ�I_�r}@O��A��
\V;���}�F�st�R��q��u�6���6����Ľ����ɏ�h?Mփs��p��/1� J�H�8���%Rəf�)��货1��o�C�����"+C�#����7�Q��;�2v+�C���p`4��eWgR<�`eĨ�#�
�7�����M�z�eE`�9m�ǁv�FX���,S0�H��6�%�!G
ܽL�M!���NL7&��'Bfr�T����y�)�^Q�׀��/�:8G��K߫�N>S���7�T�cL�R�gSs��5����_��+k�p�ڱ"����T0Q� ,����o�_J2����D�v�+��8d����kl�$�3ᦷ:�a��Av��Ȏ���Q���9��lS#8{��U�Ph���?��a�}���>��R����J�{�TD�So�1�X	� �j yh�$+qᦐ{�_
�{JJ\���w��D�JU�d���צ��F#��f���9q�C�0r��N'ܪ4�=6�Q�W
ߑ� �����A�ѽ�:*%�0Cr�R��T�����?F��iwK�����>�m0E�1a�U���zN*CF1�%�a�k4�?ƻ'�����-��7%�퀄���-�p��w����W�^s{8�e
��R����F�=jj_�bQӐ�{����S���<�i��q*တ�M���y��o@9�D��N�����k 0��Zw ��O�q�����? ��`�O4�?څ{`���H��@�ʍ�H5A��,M��@������ǆSQ6f�D���"h)���zO��'��+���efb�	����4��G�jP\��[[�����#1]�� ���L�"]��iM-#�ߎ�&�zd����]#���=/UUH�XN����S�^��i ����pZ\}��g\c�TC��-��N�Ż$�a�vR!��>ǜ��uj�+��.�7��ωlيd��Jz'�0��4������p
���x뭷��8� ��22�k�@	>z���}��+���2V�X�`���Y���|(�{�Һ`:g�=���#�5,T����4V��%�6��0�V�n�sH�_I@,�9�n�?v���j�~��#�3��W�q��`���qv�Q��\v�N�M1����U� 8g*v݁��ߕ7�	�*��ft�^4˾Ac|����������J�y:�;���\i�l����s:� e���f�#ڋ�B��Z�-ٙ��y _.��CSQKX�TB�ٝñ��O�����j��;uD�͜L@�# �h_��=¢f\CY�"�2φ�D)@�O@k�-w�<�Ǌ�D�=?c�O0$�Ta8M��o_J�|L:�@����O�h���}��m-�9��d�k�%�c�C4<� J�c(!/w$܅�8't�Dű���W�y�i<j`PB�q�f[�H`�����8��(B�2��ޱ%%��Y��H�����	t�>.�y�&���]?�<*��Bl�=#8�-kP_�#~�B� ���-v�>��*�W����m/�Ι��r�"�/�g=� mN��Q�cš�N�lXn�Y]`�ʽ��2y�F�R��"i����H�1p"Qp������V����ԙ�Vط�Z�i�[��+�eo��Qɸ>s�Nި�� ��*YaN�>1,�
�=� <6裘9���e�%���@�^S?)�QĶ#Y�1����?��=���x?��\{���!�ߍP��+�c�%ϵ*��{"�կy(KÊ�ڣ�UH�`��S�3�{�����f��M혧J\cf����hf}r�;���ptHMWg��sXw0��ܢ�ig�4�Il�Wrx���f��X����ۚc7�h��w�����Us�,Ϩ�^�I��J*��y�'���@ �Nё���Y_���e+?؟8:xƞ�Ϊ��ײώ;!���m3�f�3uo�-�l^�6�������fSI��F=�UH�`�1p��fy0�4)�pt~�z�k'n���J��R\�=�)$|+8�o���͗���Q'b
W4�~�vYC�$���2y_���h_�X�{~�P�FI�X�!>����2�>�+^�|W�/5>�M#�����Sۚц���}��Mqfk��~ÛX�X��Ԅ8GO��O�BE�ű$}?���x�����a*2��LS33گ^.�D�{��EA����:c9������޼���U��Yv����v��0���	�r�c1H:��&w�AXi~���f�I�E�0�E��^�����e�R饆�W8T�R�K,��#eLn��,�s�)���!��
*�3�·M�n�ګ5r�����ʠdM<n
^��Q�R�����4ӑ�(�w�}���q(ݤ|�P�ҶF)Ǜ1��]�3�gO*82^8B��f*9q6�����x��*��Yƅ�BG�xw[W�T+�Ym��r������¹M�4.H<EȈ�Il��z6+��տ��5hl,#�;g���\!��S�_�T�d�ɹ4��t�pp��Y�:��@��+U�>�@������Y>!ٓ�"�g��D{pbE�(9��yKH�\�x�u�@��Ą�1�̮R�M��t��yXj�.��}��'j�i࠮��.<xLrN�T|��9\�(��0��w�[y(�!���ʬ�J:��:�l�t�iE~_����$��a�,vl%�h+��	��>[>K�n%!��#��ѳ��#< ��q�z/; ա�w���W�댐L�f=�(y�F�܍�"��r� ͹�0x��̱�w�.���p�#q���r����SD�4���`O�8�ݝ'{v�\���D\�}63j�bk]�y4��� ��+z�Ļ||�,I�����a�!EY%	����dzRg���M�8A��޺`iJE.�=l��r�E]@>��W�Dy�~��0n��Mm�X�|�x��+�QqjS����m�nly�q��߿�a&$wH%�$Q֟~��W�|�*��BNL�����|Z�%	�� �( �AX҆�!�����iQP����G�ˤ��)��(v���'�I�����\�}�������L�9썞`�[,��z���x�ϣ�C�����\�0�q�&t����BQ�e�9��Z}�s���R�i��؃Q�t�� D������m��������D�"��zY�ɜC©Lw�$3�W;P��;��)�5�����MH���#4���:�)�A,�����w�.���1؁���Δ?�J�vm�C��t����]c��"��8��JEՐAl)�n�Sڿ8�B�Ѷ]zL�E	-c?x���z,�x�*��I��XB`�$屩=�uE�|�����[��0���ͥ0-��
K�{��u��N���S=j~�I�s��]S)p�{��`ݔ��H���U[F�!�`'~,�O4�zt�{��;���˔�ݨ��;<hX�v8�����Vڟ��sZ�q��ˢ��'P
.g�q�|VBr�[�7�*�jr�4wX2���
�iV�T�Y2��#\��{l=KCB]���&�C�/���,�8J�~-{Od�z�KV�Qȥ���*��)��ĥ��6P���U��\<����C(�L��-������Xřc>Y�����BV�Y���K2?�b˴��������o���|g�^5�*�81��W2j�Y��@S'wt���"���~"�5wͬV�t'
�R�&�t�l�	(>��C@�M�>�у��)��w
�O�8ĐZ��rx�n��.���[�����9*���3Wg0�!&����� a:���K�e�n٘�l<J�.Jx^U�6�$�/�G��ɲ�����W��2������"Q��ZX�=�I��z�'�Y�B>�	N�(�8X.)Aq4�ly�N� '���rF�^�=�j 8���"z+���(�iΐ�k���qS��v�l4N�6����=W�T�-3LV
q�@Y�p7�ҡ�j�wxFbw��q0I�I�y��o�+��6�5��(���d���mL�6S�c�O�F�����W�ک	�n��o�}�y!��+�����?��u�?{y\,�ҡ0�"����`#�0�&:*gSp9�8���}nIH���U6?.%6jK�����`�.�[V"&�O�2D;P��,Z�_9�#������<��q��P$��j���kd��<���i��F�����g���}m��Q/V�i��{V�.����f X��!�2%u�u�͒��7�������V���Hm �H�9��'���8vM�iB��In(���S�P�~�ϧJoQLsx���������o);i^nH^6Rj�W%��Ert�-���v|I��V��a3m)կ[� �o�0�)�ֻ�2�4O	<i/hх���b���>���#�����j���*9�������N9}U:�5�V+:)U���+|q�������l{�	�4[/���wwpL��<��M��x�V� ́D�S��f�<!�J�qJ��"��,;��n��:�ׅw1�y7[<R-�`�Y�G���)�E	O��4�욺�h�B�Z��,A��
�3u�e��Û�8(������Y4n��A+,?;�zj���k,{��J%��7rU4���f���q@�J0�z���������TrMZ���A��stߛR!�-��,|����\��'R�w�C�_Λ�U��Qy�����rZ��5r�ȧ^[���/��<��\,#<I(�(�z�Y�ܒ�9�cL���s	���ń�?���L�A��F��P�L`�Wҗv&M�n�xc��BA��)$��~ "zS[��� l-5��p�����v.*�B����?�L�6�&C����䛭J��Ȏ��?�kg��w,�$��Z���L�HMS��ʾ�p���	,�����7>3�i�<E�(�ɞp��p[]T+[�ޔv��<؀=P'��{)z�:��ap�>���B�� xLU�9��n��9�(��P���0�5&�~i����9��E��u�/a�\"��=u���{�]O��L��{�K4�� @��߶ߌ}��Po���"�D��*-�ctl4���nf1�G�̦�M�լ��ΆC�S`U�#�J�$�f���xR��k�nNPbD���6S���%����9�YZ%Q���Q�`��z�o��A���/�"�f�D^����K�O�K.��6�#,ڒ�P��""���J??�ܔ��1�=��m�?;�n�ԙ��:�=��9�	�f�W��+�n��S �m�\?{h�1�d�*��Q�H��B��k�s23�%:��T�Դ��u������}�xV�V�WBCv<8w��]?tʹ�Q6/�Z0Ӛ��Ņ�vO�C�W�W�&W��*�L��9��Fu�2fR���T��dpC6�olM?Ӌ��'���5�^���u��E���՜H���Z�)imљQ)pCd4;h5OV�
��M�@m44������#(V J�εۜy=�Į�ѿz�(���R��m�
41(A�.ͻ3;�Ǻi�(�E#5=Sb'�+�u/�9�77H�ִ�,`FXWҜ\	T�*`L�R�H��^ ���j#���:V��U�Ć��+Zq$�����A���ߕ�z���d���g(��{��RG�UE�f/�Z��IE��:~�?�~����;8�Y��ic��Zb}�P�6��p4����X�F/#"-(��@��M��]Ko�H&�w�%&6��"2���ęEfʬ$�t����!�c�_޾;�]���C��&�7�Q�$z��q
�9�xvf�>7M1����ea$jj~<�	���{󚑬𛪼\o?�:��K��H�Wiqfd��΃A���a8����;s�no)�{Ke�n��f��X���kz��頫�w��C.���6��Z#+j?�����y�0��KK��DVC[ǡ�n��I���s���{��s���ib�H��WT������A�jܡT���sWt��-5��)��jj��C/y�Iw�����:�Y�:��>6n7�Y�$���z!���	~��7kq`�:��FJ�����zď6�h7��..4.�2�����߯}lϰ��m�1D�Z�H_U�D�"A����^�����Af���������D55��/v��$z&X�B�(ȴGϑ�D������]���}�U��Bi���|�6�&�B>� �t7~�z��8�`��Yw0�Ec9�!0'�i��W�ӑvF�*aH^&�ҁ��}9�h��
`{=��&�y*H�J�&��à�?����z2�'�$�<�1m�H�63g$[}H�Tt$�*��\�[v�!��A�]DOA$��U%�� h�<�Z����X���*�5<�������}w������ �� ���]��
�aM�\?#[:�TҒ&�"�	?�gՅ�pA�.�MQ���U���4��՛�oj�0`&$[�$ѳُQ\�3�yY0�NWGX)4��df�X�u�cKy����X��d�k��@�.�o4�9��"Z�ϸ�ƾ�������nei aP�(k�N�h)���=s[��,4���3,r�n""{`��k�G����=�06��Q�ݹ����Ni��lZ�vH�r�7�Ib1LV`"��+��KB�c�&�cOk����+�i$������Xb�������Twj�*��׬v�C�V�&���u��6,�WA�a�ʛc���Γ�<��p廑���Qʣ�ed���C����4dF�?n����M��� n��!�R�zt1O?�.i��xb����^zN���#��NRX��ҋ�ۄ�~Ig
���qwY���q�.�mJf��-����6�U�1���ˆcf��,e�NM�_!	��zc�YDI�t9<�Z�V4&���kHH�beFX��A,=���].��)�E�;�]�)ǦW\�fzZ��uWj\{���I#���FV��P���BMy�RD&���(���zk�[R5�wڀ����՜s�
aJ����J�� R~P>_�M������]����D:��c{�X�<Pe�i�{�v���~��	���)a�ȓUd�Հ1�kqz O?H:+���� x�%��4����ҭ|�"����ay�x��=7NKZ���:��b�܋r���aZ�axo@Ǵ�HY�oXV�������g���|��i��w��A_R����ڴC"o�U����t]��k��F�*�_>zPj���vRsu]?�W {��`ܵt�.�jf�^�#���7fh|ς��rWN�>p�)߱F7�fm��D{3�~{�T�e,A4�ֲ���e od�+��|���d�nm�#z��v��3�
6��@�La�����9eę��ۭo��(Z��㓓���|��
��ͤ�gc{I�'�Ԩ{���'M�!?�[q2�7�﬛�m�/lQv�nt���ڒ5�9� ̲�q�Cok���W�I_D�J�,|���Zה��@Ci?㯏��O�k]�v�lP�R[%�l!r2�,*�x�J�2��Þl"҂A���V��3���5�z��^w�;(�xА0n��"���,̨��69r�]#d�'�+�i�BȨk�K�M�A�C;A�+AF�@q��j�%�iyu}�����O���xӝoSEKب]2k=���l$�q����>��_��2�D���3`����[�,Pb����&)�gU9��c��z,hQ��6ky�;u��c�PI_ö��%?~U]�X��9��J$�����x���kcr��2Uꭞ�� ����M�P�����LñN���J�/A����tW��/��Cs�r����m��۾��]����̀H��K��8�}�t���L�
��U+�p��E�0]��D�'�- �{xK�[����[
�7-OD<d%����9Y'&v�G�%=��v�:�KkD^�� ���K�Z��u��ܒz��䏦���H�����nb�c�L�=����1Pa���Dg�GV�.�2�iCe���y2����' ��W���a���&�L���-p!�9�;�%�OB	
��$Ԝ�srW���̀�S\#�X�+���dy>z�l #g~+��q1�m)���i�Y��$S!^#%\WI� ��|�lz i�4��rEd��V2��{Ŏ}]�5ތ�}7HS����S�y?��7�u��4���9p�`��Yp�㕏g��3	E�[m�I1h�
�3J��(Y�갃�^})L�s�I�Up��f�r�tR�`�-.��~&��}�W��MZ;�4+|����y�Њ�\ 5�N;{x��e4�
�4	��t��;}X�eP�z���n

xk��M��x���' .ƚ,�+]�E@���$g)�REPJj*qs�0�ʁt��ck�VL뚭#D��/�V��;)K�����_Agà�x����Z��E�8���' t��L�/Ԙ�m6n��m0��&j��9ly���@oj���&���N�3��x'˘��/.�-H�F��?LG��=ӼL�g���3k����La��S�W'.k@��L�t��aq�Ffy�$F�U�O��[7%�:��j�b���g�l�VH��p/䴢�b.�T6;���D9^�bvX�/V��쬽�ӗ�roc��ʬ�7T�tY(��jP�D�j��M�Ծ�?����] �=�X;���:O��Y6b��?kG[�sX���R�FI����\�!0
���{Zdq����W����~�F�Ŕ����r�^Ԕ��cò#d6��km����9�3E�~Ut"H��~�D��$w�vA�ͽY��
�m�g;Vݹ ��;�MI���'?�RR��Q�NM�R�-�q�rB4�d��}�f5w��Fºu�9�MᐍY������z잔�hy�i3��V�/���e8*RF�^*��/u�S�7a�`�(`de���W]U���7��'���K-#iq�1o�q�]��������b�b8��[��!�;evf���i	���1���L�$}��H~�#�9nII��F�fw��ʳ�QG�!�h&�;�{GZ��a}��N�Ǣ^3�">�'^���AE��������!`AE��^����sx&�W�j-����:	i��J�Y��]ś�v=�ʃ��M7sR=4+��)g��<^9/m��� �� R(��R	�t�y>�6A\|f�=.:��#���6�q��A#>���Y8�GH>
7/*t��ϼX̖����+7Mt�l9N�^dvL����'�>��w������{pe���$��qܾG��;F~$�n͍�L�D�O��E6vl�{v�+���{c��g��a;,��6��L��}I�j�6I�6!:M3���w�`���$��z �eߏ>S�z	I�=�p(�'�gU�6�<)z�%�4�)@|N(L�mB׊� t/u��� R��>�2@lަP|CF����*q �~��1x��)�t�"�Y劳�p8,�����G�l��a:���g�p����{𭬕�U��w��m�j��#���%}������rxV���i.�r�%���~tQ��X�yQ�V�|���)������ت���Cw�6��,H�.X�O��w���n��zK~��M���v�LV^�e_�z��Mqdl��E�>��srjHr0�*���s�w&
�"��e"�HQ���&����׫�+�����k�2��_��<&g����RT��&e�!L��Ζ�2� ���<���P��:�[ ��;�^L!�"TȮ=��9�	 ��v ���Lh�o}�<���~h(���G�xy�]ڊ4�D惯�|)Fg�OC���ǿ�%��{�Á��!�V���8���fS�E�HT5Z���{8Д�H��7zp�o;��-�����E4�X�\B�+�,��T��rj�oFg�g���7�w�YP����RV�?��P�Ч꺕d�2����>z�S�:�,�/-�,	h�|�|M靆:���/n��c4����*F�x���[��T*�C�bz�;n�����T�Qa'I�\�aa!�Dא������;��6�A�"��hĀ���0_6�	�Sb�@3SH7<*j]�,�V?���_���'RT�C����58C9����Nc��Y<�U()��"�������|*Aч�9��U3�v�v5���"�Չ��V���a��V2�ei ������(qs*B^�3[2e�A��-�n]+\�7{eVs<ctt�T=c��څ��#~Ц�|Ϡ)��ɁA+�_2�䁼'���S��!ԫ(i@���-�Qe�/{��[���f,;�%��&r�a/輍��O����A�:��[㺚*M��Ɏ�P�֬5�3���]Oh�]Y�lt� 0����? �tg����}|_T�H�� �~���M��ɩ�. RO��J	��1b����3�5�ҖZ��i�Z�f.���j]�Y�z	kG��~7�8�9�lt�q�Q���c�V������i��|����a���ɵ���#�q���I�A+��lg'�#��;���n'�)�����(8=J��j�M����7j�9t���A�M|����NY/�A��c�ZQح|����cO}T�G��&��L
�{T�%b�;��	��)�d
�$�j B�"��*�ax �
r�j~W��w�W� s��^�L5�^(���x/:w~k@�i�6�0ܢ��yZ�u�6�Ֆ��tΛ��c�\�u���p%m��� 5g���O�z��0!|�]>����W��*�mH�����jǜS*D0�YC�`��_�zug�#<���"<��ҟ�?᢫ȇ�^h�4�Dg�ȟ�m��#�=�Ǉ! &j�
�?�+sV�9�%Zc�}5�ٮo��&_W�q���Woƍ�$�WB�a'�*Q�=���b�B^W`=��.�T���`��r`�V1~7���lw��o�$QY4"R���?�ﲛ� )�&����.�c,\'�#��0]E��ő!�]�yL��=�K4A��ֲ�E��K���+�N<
e��FB��h;�_���6d�%C��W#֒��t�z��v��O�.K�1��Q+�`ȕ~��"�=h��#i��S�iN�"G��h�(.���L�ﯠ���=�`�!�����&`�c�^��ßK�Xƺ�%��j�+(��V'9��Wv?�	ߌɎ��$��x0W�2��j��w��y=�,?����:�^�Wy Au"�B��~ ��򗳩�v?�v�O�*�4
М�{� 3h���ʹ�)M��Ţɷf�2ƨ�YWl�Ym=�f3�;���2�e������P���۟��O�[5�'[n��i_7�ᑒ+c�S��r��"�$�w���]�r�_6�j|2�y4

�"t�rX��&�v�����a�eh�r�����ߥ��u�y�є�jٷ���̷��nerP�jV�u�:�*���U�A����K��L����׫�|�	�*�,�7��"�>����s���؀�:�#;VY2y��>Τ���� �>��V��軻�qd���x���}O0�pd�����P`�cT�&��_0W4��5i�&�|�k�z��jXY'�xD0���h��1Y��O|�rJ q�)\-��|3��˳�`�f+���/ŻR�R�v^M3'Ү�ךFn���;��G_�.�P���Ow�@>��ƀ�����̪���{<�P�r�:��LPXNl&"�]��2�w�G��CΪ�^�y�ykKz����#���+���V���T�����F��ۋmM�6�j8+[�k��ul8|P ��Bz)��}�֧�#~������f�
Rc(3��R�"?F�uj�þ�8���ϩ4��v�M%%�٨`����N�۔O�T��]h��j*��m��ť o!�]�X�9R��L��)�˕Tӗ�]�|2�')���W�d���/I�������ҖcH��{]F��Ǡޅw{�)/ӳe8]��牨��SX�Ā-�K�^��F��_(�ٙöu����j��) ��6����5�����$���DsE<½��f�W(U=���2�w�(@>�t&Π3�;�R�D��N	�vg$��t΢P���3A�zA��8N���7�V�D<��-2�n��U����<L:w΃w}"�G�!�s�o5���+����O��$�Jq?~kԶ��y=���6�)����"���ӝW%�w��8ۦ��onY�����DΈ��4,�.rЪeo,;6y����e.��`�`s���*%�a>��Z6�)��u���rJ'��Y��cKV$��̑׿��?%@����,�^!F�[b�S�e�|T�	����ԃ%zY���	�瘴���X�V�Tձw����7Rk���2��&ŗ!�	d��n��|�=K�tQ�{F�Ռk =��e8�t�G�?����R]��� �A� xX3k3�\Hb��F�6'�o�r�" �����u5'C��w!�eu'�`#�j�bJ(ɗ�����~�WP�$�F�{��4��U�D�BC��TIT����Dh]��5��M*RQ�<D�UC�]]��t�<�t6� �N�YA�E��xB�	ﶴ�r��I9��[}k��H�5�4�Yw�c��{�M&�ͤ��NK�5�2ԫ�͡�!e)����P��O�ޒ�e�-��s�-���$a�O�F�H(��UV�(�>3Fh�s�Gv�.T+}����WB7���-c�Ɔ�7�ֿ`0���G��W��zS�4�֗�MxH�VH�*'���j�������2���	�La���ˋf|�V�d��$��Jq��C��vt9��D����V��l<�\K��P��ޚ�<���'�&�^�V���RRB*"4�DO��n0��p��,���p�#�f1���+�Z�!ç��9�0I�#����`�,�U��z���&��������[-�4"e��2%#�z����v�5�U���+��\���ج%/_�Ou�M������z���Syc�0u|�L�n��|�[�����E���m��T�ї���	pmez�==�Z�]��/S������%�ԧ�-��5{�Տ�c�I;h��l�)�$S����xrP��Vּ/����=�\ �۵����5���B1�r�M�(�O�PHN�lc�4:a��[� Hav�I��s�Y�D�Z�/ �G�]*�-亟*	ހ��ܛ�0(g]�].ڋ	�P��ktk��S���=�3�ֱ�(�"i�!���I/쫺?��1e!
j��2��0sR�L�̫�����*�W���Z�Vuz���L\ĩ�u;�}wTGB8�)�S���g�S��gK�w��66<9$�5 �(�sBf�Q����X�%����~7O��\��!qڋ�D�3�e3595�dF��
���"h�=I;�)4���A�@�z�[;��~/:�&�����*8�>y=���z�/';�efp&��A��ʫ�����qcTG�VK���0��!~��g8�/�+!ɲ�0���i����ُ�]E���JqѸ�NNP[k����3G	ެd�V�Z>��4�?	�����ธ=l��!���D����޾�ߊ�:ő�h����d}:���/�1kى�������z��6�`=;���v�r�\�Iܥ4�JUq�eb��4q�	�$45Y�������A��#�U8U��5a��~G��A�~�"H7�	�Ш뼠�5� ���]�Tje�m3��3?��R�ؠ��;��� ��c3Ʋ��A��aq�s�ع�~+~a�	�J��u�sE�iP���v@i�B�X��L�'���&�� �>������>�`k�=B�I���*��d�������ˉS��^��
�z.�W!�+T*�Z��^��`z�=��ȆE��0.�~�:�� ��KZI�r(�<E:|p>�)��C�Q�x�q���݁�XP�n����td�v�K����ٍT�9�:~�>��b���D�+��<S�ꏭ��оE�2�\Q_�hq�{���s�t���d	�7 ���=�x�D��<3)�/�9���z����Hmy����5h��=�@�xњ��w�H�6byOYkM�'��@�/���}P�L���X�R��5	����y����x�������&��c�]b52ޓ������1�08 �7�ȌZO���C�H7�zJY�����u��58��/���1�E�ɓS�ľ,����$�?��n׫ypj�O3y�����(�ZW'*x��/s�ߓ�"�� �PV����a��D�Q�Vп����7�]�`"��J�Q����$��{�i�����d1����@h1�A�2
r6�,������c��Mf�4Z����2�qx'xC��n�(L���(�����ے�|J�o69o��2���\d(d�+#R����nD,��7V�e���~�2�kuI��4�_�^���3[������wxb�[�ܴo�Έ	ϵ��U1�H��"5#�'K��F]QF�����-3d�ֳo?��Ë��?Q���Y��xL+ �HВhO8����ܠ}r��BG�t��35��@�u^G��&Li���.W*eE��� ��L0]�L�w�����-ِx�;���eP���9�v<�k�9�l���[~�M|ƕc��"c��$��9���Xd��E�V��>!hd$.[QH@\���t���xG���@�Z�*��1��e2pi1�9�p�q� �0�Qe+�\{;>���LNLN6���Q��s�`B9��O��a���E��2y�X��;�/��%B�%%�*ܐ�FE����(ƈ4�RGs�w5�Qs�M��g�]��٪��,ߩ�]ăʺGb�~��&�ҏ�KN�1�D�C�jt���=`^q�����o@r|ĶC�N�?��lo#bG�{�#�-��Ugg�nu
t�������)&�$��20��s��I�"+�y>�.:�r�1��WJ�l�G%�H��<ɘ{��\�ꄜ���W�?+��j>�P��Ϣ�����L�i��{�s%��������A�QX�
54� �[�(�&�73�
t�,�k���K�����;����j)���%_��K�����r�:�&��дoFF�(��>c6�*#:�u��
��)>��i��:@E�nb����i^�?#Ȃ�#�JK,ªj�S�&�v��^�}i��U�� �.���j��ai#��OI	eݧ�\���,\:|����"H	�����ôQj���f��q8#�T�'�}C���c:�Rl�ДozS� ���j��F�b����za�)�,��x�> �f����Q�Q8	J�^��6�u`��}���KJ�5���~�؎a�3���Yٰ'�b�{�fઢ�pl|���-�`Ctb���]{�EH<�>�+Z뎊�,��@;PL�ܐ4&��$Q�}�k��8"P���WOt� �Y���k��U.����mJ��L�6���� =�'N��җrq1s�ݕD� �=�(�xzI��dD�e�|�3�?-,�3Ɋ禦���f1��%�AD	�d�&�;��f:ڬ�˂��U	(��K�fG؁4-[RVu��} m�^U�H�% �<�/��3�UMrUj|b1 �߽i;�,b�59LnF�V�~�"�=����S9s���Y��@������Ed!�	��<�͸����i���5�T-�ݒ9/tՈ6G^\[�� ���g�k�D��7�;�z�~�ԡ��}D��a?l�h���x+�M����s�r;ړH�#-��	�@d���;l��
���"���U�S���`�gp��j��[?����P�\iIV��G�2]-l��]ߦ��#"Ƈ?[����\�����dc��-�l��Ɩ{��,��m�)<�l��JX�@֡�9�aݥ*�l��s;M���3l�9��[���v�O-'��^J��:�H	�!�|ݳ�ޘE����s�fK�h��&�I�i�e�M�f�K�P��� 2ݿE�� w6�����l�:=�������ߙ�t���7���0��4�������v<ݖ�^*i����������w��nN�H�����+�׫,/���Q���r!ٟd@�>v���t��P��p@�P��,�])�Y;O�Ţ)|�'g�/q�,���yM	�h/�씐T 6�--��2��t}�{���(�����p�pL�w �InL8+;���s��1^�7��ˏ��r�	���4t��	y_M���Gkc��Me�r+�~�Y�闛Wd�ޖ��Ļ� ���k�g��eX��&+��ye{P��Z�4�Q$=B�v�@���^��"�ui����t�<�m��zޮ�|o�mէ�/���n߈u7C?�/�6�$�[Հ3��8��:���|�й�ҫ�\�m�b7KZ�K��<(��P�fp�/��q�S��O&�>ZHz�_>�p�j͸��u
���k�n����O��m�7P~�����Fw�z���ܧO'g����mť����<��k��������[1��L�q��ũ0=E:<�z�}Ӓ�-%�2����o{�g�.� ��-3G�P��%�P���|3(
ŇU��&�9����w� ɛ8��U�2���Ɯl��C;/T���#�/�.�-���E*�:(��)��'1·���2=6�T5���$����fjb�dPU'�M�<���?�T'X<��I��r�d�lB�>q[��
4�&x:@(G5����i�����I�Jk�x���F�����񈮸iKL�m�#�H^��>Y�u�<��u���Z�5o����RO��ح���h�z�E }ϼT����J���^����%?���Ǎe��č���D��5�ipp��b~��Ԟ��3?��J�tߋ��!u����N�, ��ʃض��d����G���3"He��(\��)E)ls_�9JΠz|:#Y���m��[�N�����F#t5FGS�p���N_��P[xP�w�.=[�I�2�J��ᑨ�vH�3!kyX�r���!.G�58�	�-1����D�^?Z\�Q�m�[|wc5랾\� 6��m�����/�e󢒜�BLB�p�mHA�+w�nۅ��\�M����݄f� MEO��`�C���!�t��ڲ*5-Gu_ �WN#�U��DX�+S$.�A�ۻ�+�� ��G=��&�_�VT����J�xr�m��Ǭw�E���p����7(Ⱦ��Đ�O�g�,>�;��� -��q�$~����П�C#�Q�hG2�2BCV
ƩȈ#��j�6�3�4)5����ZxVJ��'<�XgS��6��^Z;ބ�&�2����rK�z�>;�Ts�v�x�(-M)�K��qZ
� ��=v@�q��tV���]�	�0���B؁Q��ܳ�D�Q�o;�b�_x�'J��ה���H�>k���vkD�6�A�J�H�!�y��g����[q�7$$F�z�t����"2VR��,g1E���.��!�
�V@�Ȯ[��Ć����*k��G=�o��H��Of�Nղј��mS0�z�<�Z����b�|�|<��������EE�"ᩆ?�,��y��u� �`��t�v���ER&���}C�t�_��X��:D�KUgnM̣��r�l���F��Q18�d�\4t���7D��XS�x83+�8m�]y�e�g8R���(��x��S����u.I�r)���t���'����r�m��0�-Z���P/�����M��L�h�{�i�~K	�f���D^��]L���F��ɦjiSXZk�c��]�Z�~�[��&1G'���0/
ȡlXH��f�_F�cMC�W���{2����?�j�z�`N��Sd������mp�S�М����n�q~�о�+b�}&��}�.�������#�⚷����}-�Z<^�����.n���b�liEy��+�x���ތi�A��`�`�����<}rw��SV�N�1�!���Y����C�H'�AI@B��-�q ��'� �Ej�SY ���,*әL.&��y!Bo�l��E�����TJ�Z�(w���s�Zam��k�*���4����Ѭ��6��6���-��_Wp�N)�v5�p�<��aNt��"�ԏd�p�./��	��ϣES���Y��r�b̚n�f����)�2�_?O�%	{lDǓp�ya�X[���ga׌�7M�ӹ�<eI��0�d% ^��_�R,@�]Z��4}�ȝINUϭ�քopy�3�)_�v�e�(�=}��1��qЃت$*��"
R��[86L�l�T�w�������H
���9٘Z����6�RŚ�ɰ~��8��[77��+�p@[�EL����JHI�8���~T;�=ɡ0�����7�"�Ӕz+,j��O�+n��dM��zx���a�v�	b\',�0������ץ.:��a.-���m	��e*�2u~x�S*=�M�I8��T���9RHx��x�x5g�N��C'�Jo�P?�k���'C[Ru�G�5\7�Z<&[�qφ���;-=�T�*a�83/=����G�s��½�=~Z��ź��]w���=��Pojrh苤�	���v,~��Ɵ�K�f,�W��j�W�ԞA6I���<����i�u�RstzS`�& Q����85�J �9)�Q ��V;���+G9�g�%��Y������^ǒ��TU@�.����[49�Փ���t��	9��ߑLHo�/����!E�}[�0��O�ZXI���)�<Ո?�޺�y�)���;�����K��t�E:ӸJRnZ=(�#b�[��'�����	�)��u�o�{m"{��cv��d1�9ָ�S"��@��R��0q��^2O�K ̵)>�6������=�������h;~��xA�=���)�T3J�LBm�e9{��';c\����:f��X�~��Lp�ǅ˚�.̇�×!$���\��I�	�a��\3�saٱ���-'9OY����P�%���ux�R(ib[���Bê�T�,Ol�Ea ����Fe��[�#��,���Aˋ� 5��\��v����N#v��`���xF���1]Ɵ��;�� �V����w��f
����hB����Ӓ���,��=a%��6N���{F"��G��Kes�SMÝJ���ce���4~t�LrYk������^v��K?�R������;��У{��m,��ѯ�������t0=?wǂ�Ch��E�,��	�e���C�I�=X�hgo��}���BÍk�!�#d�%Ar7$"?���#q E��ЮK`�[�7����wX��$�ph���,��n�z6,��j�*0h�9���"Fa$��0(�i��:Z
��4����������#?n�qp���N�.=���� ����i��g���V\�3T�E��:{y�NCJ�7������5�@�}2��5�M�Rӊd(ک��zO���������{��Ғ��Ua�T�a����sșF�|�S�d�,v=�1����BbE&�Ʇ���������k*r�x�j
F2�����Q��k`���+nZ��ń�Z��Q��CGc��ŭ�Z��s7��6�1.=B��_AԲ8�|rH����@���A �f�1x�����ߍ��������S��O��u����V�&,烘B�&�� ӵ��hKKJ��R��,UZ�C�d R�.e�3��8�e��pwtp�W��h��V����@�ퟻ�kQwz�YѶQq�h.��������O�x�a�]/Cu��.��0�iS�NR/���}Q�b@��"�2~!+)�H�.CtU�s�@�0�N��iPZ(Z��f\�1m\����M��W��c�2ku�D&[�������Y��@1f�H����wL�"Wt�z���ΝKC�Q��[�����n�o�J�T�_4@�5�+<K<��ɿ��x���1�'�����֑a� <�>�	f!Ԗ=U�%g��x����p�6c��bml��+8>(��3��e���QZ\����,ܦlp�[��0v�z�9��[�����������h�R�;��Y�Z�y�%�a*-��A��-���j�1�0�oZCY+���K���8!;��cmFp,t�VX�,�iA�MS?v�:���������oo�����C�o���R/Ȯ*6��5�3���ս�r=���j.� &�|�aZ5Uag������7�ի�MϦ�ʖ��u�6�gK��[��̯�_,~i7A�x�_�9����;�5�mȍ�X2:����Z�TZ��`!�r�Gǎ�N��?l���%�M �Oޭ�>(���7�b�'J���(Bֱ��b��ͽ�3���a�ɐ���h-�c�#1��t>rpLs��BI�̕�ց�ϛ�Cj,�h��H���~g�/�� t�R/��) �����K?�o(�x�{�ls�G�a�GTs|<^e�We>�ɱ��	r���o	s�F"�-�yE$}��{;f
�{�S���=WVҨ*��q8�FsrN���v�K�bq�P5	�\����b�^2�ڌ-��]S )�_3(��ߐՌ&�8�1!{�f� 囧�)�9�o������v���r �����\1�e�Vc��Y6����E�T����t�=��+��Y 28�b	��ћ�.1.��߉6ܔD��E҄ϡ�����ik�P:R����5�ޫ0Mp�m�q��ؒRL�d�-�RO;}������&:5s�&p-�B�0�)�؉;ѷ�O/.�g��1��)���C~R�r��N�qt0A/)ը'5����j��lQJ=�^KG7T	���Щ�0�=謥�K?��w"�/�*�������q�Tu��h��ppo�jcp��S��m��?�c�>�ٙک�:)XT�l��q?2�T����&��������xAM~��
;���N�OqJ^�����w��L/��4��RF�%2>K	فO�9�/�ᥠz�Wb�X��QK�^����>���eݚq�\O��jz����He\r���sb�����-Ř���F�������IH��>;n�����7�կ)��X�(#�4�sbg��(�ΫM��t,�˛���蟗��U���싾V7��\�e=a�|��\�P�]���v�.�4A*糄
�ЯYS�丛8�dF=٦[K>\�i�7w0?|��D�����+b�p���ӄ��ձ��U����k��(���oӱ<�䠁�M���&y������当S�����A!�ɬ!o&^�kd����1>_ �y�	��]�)^1Ʉ��I�<��P���*�R\��x�;�HX��_��.l�ܶ+d�-�9�Sa��Y��ȱ�g�W�w�����,i"���-��BFvt��^3����g��@I�-�d�(�W�{QU�-=`t����I	�s��z�Es=��I�����ak�>���Ҧ0�I���#�Ņ -�1���6��Ö�ʻJ��n����n��m�ރ�3���8��6�T�c_@x�p{�Fʽ�U���͉x<2><'Q���g�����#��6�p��-it��F@�Ξ�qizn��7��cA��q�@L�Y	0���q��4K}��q���Z��0K�o*����g&���x�@،����[v@�9E�Ą�����O��uS]�%b�
jhY���f��?G�����5?u<"3�r�R�H:od�,b@A]����[��Ը��c�IE�G/fe����T܎\�[t�mz�����/ى	��m�?�}���8E!,cz �w�3>"����M��E[D�U8�14y�8)��b�>l5�ɂ�r��R-�ԁ�J	g���bߟ���ڿV���Ȓ��jic�@��}��o�ǆ�6�1;M'�q;=����'�-%:ʢ�T�A���m��$�<U	5�,����ھ~�}d���P]Gm�"G���Ͱ�b˒·0�n�Ď�f]��q5Ӝ��^
����iL=�����b_�3�%�#g�fz�F�S����(3o\�,�O��.v�A�f�w�z�r�J_]��Q��T��b�C4�/"�c��2�E����m�l���D�0�3E��L�斒�2��>��A�QL�1NDT��χS�"�QC�r?5aXx�MY3�)T��1�>���Z��>HL��)����u��H w&v?�����ܜ����n�-p����T|Y�ޯ�Cf������w�6R&��O��j��4���C�bB^�v�'�w`Fq%�cw����ѿ:t�p`ხ�pvK�@0�<{�RE�����'���b����A�,c]�!��x�Az6��H�绰B�^a]l6�KY� ��{���UmV�"�QhWS�i�>ñO0��+,�.�q63ZJ?�����q�BV���x�r)�PGR	�s�
_P?����u�>o/%^��]������H��A���r�γ��i�ɞ-�FR-���q\$Q�Wr�:���(�0"�N�{������@�b�3��F��$��]��b	5��*:Q9L�;{�(y�^+]"�sP�=�X�a$#H3���t�0�ХCj(p^����fLEŀ+���cӳhxlДV?��}((r���U.�X�[VQ�"��/�3��?v돉{2����B�|�/�!�J�sd�!�����6fo����߁A׀"aH&Z�x`��# �%A�}�� �@�Z�\�-L���/$dS8�oHV2aMw���(N��S/�,��]�_�k��s�^�];@Ш �sr�&��|@�{$�/lQ~�'���;�I����m,�d�<�Ɔ�\]��Q�gQ廔����M�uW�q�<EJ��������{�jTsde���&�GG7ؘW�O���I 4�-�P�"y A���A9��cV��l��&�Q��j40$��Ӛ��O�� ��A)��/ ��dg�}�eTX�����:r�n�%�@���G��F8a'uT�(R%��mX�D�t�a�W�@�޺"�
���-��U�����U�LՈ����8��i�7�˕(�� �&��'��ξ�O�#K�*��K>C��L0q����4�;I�[N����Pj/�VOI�M���]9f�չj�Z�,�$x���#.����j_T=u���RJL
�l�����Y�T��_��i��Cz��j��1P�����ա��%��z][~��u��x��3s�dP8'�\� <{Ơ�̀�Jb�ߨo�z��ה�^zQQ ���+�-��j��#�����B7_�C�L���<���]�3�(L0^8���w�S��zW���r?�mL��3�ݏ,�a�ڕ���d�	3˷f;0j�q�1��TD~��Z�9�����0ah~^��d�ơ��U\;&GR�x;�g)ޞ�<��	�!��� �_tO�O_��?����N��J��Hiڻ�$L
P��x�4�m�=/�,��`�J�0�?�@'�'M$�+fm���i�Jֈ���b*(��O	�gFp[���$N�c~����|��j�S��lb�5	|L�CcW�C��$��z�	�N~��V�v�?�󝅆����;S�/�nDN��^�+���I��O�F�;9*9�d���"�)A����F�8����O�T�Eິﾢ��1�-M���E���+�T��E�b�'4̲�3��c�������z[~^(���X���5��glݺ�w��=j�_V����/� β���M�����s��D�ONa
Y��~�j��LV�u�X��?c���e]��L������39!!���[�i�\�c�1����X7��C�r��%k;����@+���bYZ	Q]�ؒ���@�O��(1Ȱ;Ԕ@�ӧ.,��<ӄ��|P?~��k�<fN��g��A0ENlh�W$�/�����+��.��&��wS�	�7#��@��3ɬB��/U׏�9��$�O~�c�%Ǭ:)�U������*�����Ҝ��#X��W�T�4XG��L��d���f�+���G��yQ0؏��%_����|���Y9�`�"��HF���TIYOP�n<r�Qv� L���4�~��U��G�榚����	����c��K�
��rU�Jg�Yݪw���!�	��������ו��t���"�. �>�`,�sl=��-�tDI�W�DB�g��8�*��Q <�2*Ny2X�����-N��H잏p��^�qk̔x8GR��upf<��{б�x�v`7�\�d��=\~".�TT�f�rL���
��}�dmd��oNn��o�4n�!����d7�P�ъ��7�/���+_M�C�[~��*?��Aʞ7��⹺C8����f�
���m��iѵ��H����Y��E��U�1{�å]�6�:��ɲ����2[�� �x�5�o�$����X2[�Du���H�U0�W��:�,�TnBnr��!'|CP��
Wx����Q�d�%����l�&d�ִ��f<���c !�� ��f+���T�G���}��������
�ƥ���6�yx�9�v+��������~/�AL@��R���P��[YU=��렄Y�,"$P��.��3����hQa�S-�$wҍ^$~A�.����T�d�*-� AA���$�Q����z�Y���(ʯ���"�'I 0@�|��N5�I�ʔ���e�y��)R1O�wJ�@Ͽ0�V�� ܾv����ܾ�ĘF�۸fVB#�%Ƙ���94�`Y�AØR�#zTY/�n#9�� �O��K@�t>����K�������2f�:�����Y��-���-z9w�Vŉ��@���������o�q�֣O�S�7a���d�!Q�h��]�ks@$�/�]?H��S{��V�!�4P4����B�8ݤW�5+y��C"1��aq� 5���ks�v�c�}9_*Y�h2+wE�j���)�Gp�{�x���
��MZ���O4xĞ�qIt�t��1-��tJ�Ǔ������r�� ���^�������a��X��h���g�@�C�#���7|*z��������#c�ۘ��o�J��͉ʀ]��"��,r3��mZ�Q/�u#ΝF$����L�0�6�h�2�����N���
�aՠ�l�*����^L��1���p�T�K#��H��G�0ut	Ek��maD|о����G;:��t����g�1
�(ڢ�g������c�M7q��5�B���-� �쾵��4k{Y䏙�LA���R}�M'��.P���Q����"�sk˛�?n�]�>�xz������ b&�zK'
s�
_ڹ�����xXl,tf���k @�v��_�*�8ܥ�&�r|�&�s��x- NFX�Y�(�z�Kԏ�(��
�IB�/f�����:$>S���S�ЭM	��<+k�r%�NM����wvL����!��0�0'wNr��շ];���L�r�S�SBE��'� ���v�w�ƴ�·�l��L��N,N�͸�G����6[z�z�(d]���n��f�/����eV��X���R��Y��\t��&dyk1�A��k���}�u.
���
?�Yx��t����qhݵ�`!�,7z�
��Y�c���U�H��ͱqd��Ѫg���tb���"��TՐ+�^��l}f]U0{���ZhYח��Z)S�H�)U������}��n.8�z��M����`��>1鷳��U���I:�9���������(�w@J����ਿ|x4�j�.��|����t-T�AA١��S�V'� L S.j!�"��Odm�#	�6ȣRO���a�@�Mځl"���#�t��� �Y@L�E��Ѱ8L

�{��������z�f2�-�	����E#D�V0<&��WR��1Y����b��<��.ۀ�8��ԑr|j`��(��IS�h�y�k-<Q��f�A�fmW A��V�+x�T��&)MrI�$L�����2��vh����n%'�G���Z���{[8���xmH2�T"�T���]X��w��z)�=����ݭ���?�.q@k�V+ɹz6��\�#V�Ϛn��ߊO�Uv�@��'�)'ԋ):S~DZ��f��-
Au�HS
�3� �R�3�i�6G4.pP���T��j������zX61��nO⼦�j��#g�&>d���u�+*�����	�6��s�!�y�s��4��z�F�Zԩ
���ک&��Q�m�P���*Wi޶�Ck�E��y+d�XAu��Y^p�p8�\��(?,;����l�Rⱴ�\��v�%|�s�����1X���R=�à�sD����wA�>��^w�
>��Yo�c��j?�i�����~�R�#p�R����I]⿒��V
)wG�<�f���n�O�~��/f�b��8�K|�3甁�F���$u���������y�(|c���"�tƂ�ʹ/K�/W�M0F;e����yώeouX}���S�I��4!�5&!\iS���@C��x�}S	
k*�w!E^��I)��/���q೵�9p�e�h�0��n���'y�wݘ\�fDɗ5/�f��1�-*��X"�]�%b�y4�g�t�[ʑ��k�Ds�u6���lt�����J��z�QXTԺ�S9��E��
���=�l���w�����	��i�1;p�!���x�9L��R��A4ă��HG<䰗r���O��ʹѮ�:	�c)�4��}��	�C��ոo�w�_,&�{�ߺ�,�� �DK�g3 �l��D��f�[ȉ��X�ݨ�ֳ� }+�?��_��u	��"����,0�d��m.�G��
Ϥm����sBw��"���Z�3��p˺G�c'"���p��P^o�8v������ܮA��D"
��W���ϖ|�qP�t�j�m��M������5���`��z�`p���fh՝֦x2�ȋ��#�j6x���e8�NR����o{�7(�<�X?�Y~������}� �e�j�­z3�aZÖ:�*�E0Z{;��5z:�:��ɍ�Fd�ez��t�%��U���0؉��%@�*X�B|�M�SI�W���Q�S_+$�L�� ��MS{YU6�i�MrP����^�R�x�
V��`�l?��޸���}��c�)B]$z c�6|��ZR���*����0t[ʓdև)��h�]�RCO'����
D��?o�>����g�O�l�}���0��:�������]jO����;Q��(l�%�ɨ���Nm�P�9�`��:{�[	��� I�v'۷�un8�Qض�Rk9��6Ŏ����hDO���M��W8����N��u� �LCJp1�v��+OP2)�Υ閩��F�X^t���� ��h�)�;����g�QgV���,�����PNi �k��HD!,� i��c
��W,tp\1<�/��zT���7�����2;*�G���گ&28яpRh�n�̳EQR��Ph�*��I*!ǅF�uIy_c�)���k-<��-��F�Mg��,�'$L�J�O_^'�~��	��v��Ԕ8���`�ėJ x���Z|]����'l���&��r���K:}�O�u<�4�ի>��Ռ��Q5�R:C�UA7H�mh[d�#������vSH�))9�꟥��1����pv��pN.�=�c�5�%ɑi�N�����$�nvcu�K�#�b{��{J�
�n�G���)����8�$G������N�M�]��|�hv��/~&����s���ϮI�t��'���-�:ڦN���,�$�6�uӖnW&�Q��/���ut(j����$Q-i
�y��Bܣ���Ǝv�am�vW?44����PE9�38�d��=	4\u,Uv�R��Z�a�O!�C�}�m��L�s��g�`�M����AǴe�@#��X��0�$��Us.�R����э������G�h�JP�qݬd3�|���Z�eE �׺�J�A�<O�<E�b�p�f�{,�4�C@�QN$s=	52��/N�k���m
d��G����g��^ɢH@a/�-a9 ��\GĀ߸ՀF 6��~����7�_��5���1Y[��3�SG�m�R]Hc9��Ia��ÍI�b����8I��D������A�ZB�֎���6�;��j=j���0t���ڒ���$I|C_�V��0�=t�i��| ����Gn���9�_�fA�		)1��Ŵ�v���o���_f�[��n+�퐿R(������$�@'FM,�F�I� TczF��ڢ�`**�6Z㸸K3�#�k�u/�6�7�|v~�g���%�p�cP�B����-'�b��d����d��6��KQ�V�iV~L=;t�|��Cae:n�&� Ħ�� 1>���_�k�>�Z��?��.9�+�O��_�c�{�L����hxiN*W��%��
:�,4�T)�z�킦?��tnڜ@7qP4]��n����)�P;V��x�{L��8�W�6Ù�nWCR� �mi�h�!L�˞��js�ξ���p�,I����? �p�r�YfnhFisC3M�U�n@�w�H Wj(P����UUq;㞈�e��rPg>�P�!Es�;�R�q!�;�d�3��Ѕ-;����MzdY
خ#|��$֍8[����QH�? ��̫���D�3��m��d�4���.=tl�f��]�rXMs>��aG�K���7��O@��
q~6�ڣ,1QO �ޥ������C>�ؖ�͔D��Ȫ4ʍ���脩�-�r
��.���'�Ԗ�]�a��֮QjAc�"3�
ir3O�*����~ǄjxiN��odp������"1�x����g^g���o�;�������7�	ݵ��DpOd^��8{�	~����.�r���#]�A��)���nMT;?+��}���H+��L��q�yA�6�i�|-$�8�ӱ��_t���b��m{pGgP�Q����E&�Ve@��)Ik@!Ĺ+�.�ðQ8�J:5��ѻ^@��sGŎ>��v� �v����	����)�#�zk�Ԅ�(��i,H�},�2:�����Ʒ��8����Ky�E���Rhؗ��u����&SGwt�f$�œx�vZ�L�����A�p�T��������VɕGt��	�v�&����wy/�����aa`��� �J?��ųe��t��oX�ݎBgWʪ��Ҕ�BW��b��>z��cP��͉5.�d�<`�Ab:�h)�Di�~�s	��e�d�:����P�~J��|��'~q園����H��T��GDm=#���{��XA��ʜ�A�@_A_�,�wC�UCVK�
z�~XY^�VB�˰H�NC)�?�ES��;n3���Mu�G"Ӫ2����;d���4��UV�FTP�*{IY:w�g#ƍ�~XҖ@���M�mx����vry u�c�)�,:0��0oaˈp��mF�ɚ�ߣ�Op5�b_Ֆ�/gM$W��ˏrU���w~A��.w�v����1�N�8���Ep���(�<�vs�u�\eć�mF{�o;+����'�#8k���6���s���EzN��FƜQ!���#�T̅�q=X��8�qq3*m~��hf�f�~���gʂ=S2�qi|��	d>v����:��$���Ol����_A��1-H�5��-�,^b�
�CZ�iA���068��6�\��u=�*�F���J�*2��cH�1�	%�� �C�Q,��#h�@0�t�T��l�����s�a[�\���U)M�f�H�9�O�1�SCz/~1z+��0�my�6�Rk�m���٪��+F��&���茶�q7��x,��x�r���q���8f[��`y�>����6pw����(d�+�a��[$ԭTD�:�0�*tm	"D�(n(��V@3�AH�{*B$�����57��r�GD����_���!���\SC]t��N'a~��s���2G��n욠����m%V�kD� �T,;\� �@�B+{���0C�޵�Sے}zL.� �m���o\Gd.�B
�ֹ������:��@18�ؠ�D.!�f���#d�\��ćU�S�lW�ע������'X���r��l��T@H�;�7"��w&g��>�JivݖN�8�ʉ���ˀ��j��W�/
������v�0Z��e���/|տK��B��w{�H3(J]x��%�+Ɍ�*Mr�):����W�rW8��R{�?��#"	y�N��Hc{_!x��D_z��|��3�gC_W��4����k�~v��D�����=�y�����K������w|�m�o	��F's�h�J|��&_`-s�W�B�ZWI���uW
�ót)c:Bs9�k��Y
����A�y�k�{�#�3�D�d���^��47jU�%$$��UI��뱞�ne�eCU��Ҵ�����N1ʠ�0��Idx�S	:RU
Uz'ɴ�3�
��3Фj�䒞�9�8-�91$@���6��c;kI�!��O�\gn��4���f��Z��`��r�J�z}�7����c\i���UJҌ��a�|�Ja�],o������>��"A��D�\����.�٢,�\zJL�����z�5z;߂��Uĥn�W�BN2(5e�x���E�Α�����ZȻ�0�@��C�#�-\xwd*�<ك%ka� cF�cN�R�
��s3��$�C��2]�#oê�RE��!��� �@4K=��M����N�Q;�S8�`��m����g��-�6��i-�:�a��U�5�O�ڡ���'�~ZZ��
"��F*�Z�T����R��+z�(�R-�h��vN����8�{G9��.��Qj��=�c��i>��WBV�{���/�r��#��3F{�����"~78BF�K0�F�$��v=I������-G���n�_����n�)��j``�f5{���K�K��}�rӦ�����*-��HG��&nbѝ���r�U/�<Y���x2E�����	� �Ɏ<�@T���\4������Ivġ��eҋTхӌ.�q�!��t�;�K�yb�k�#�b��f���~�~kq���V��W-!rq�0qtNP(�sA��珎�͙�:��[�J!)��a���!����{j1<�'C�*��v_8P8Z	�E�]4���L$��[����(:�P�eG�^M3^�@��V"�ZO��"��r{7�ee
�h��B�9J�^9�7���l��9XVM�`:�5���[���Z�h6�NѠ#X+�ߊ%���N$E��)g�q^e7e�r9���rq{�F�X���}��TՑ�/���o�V�>Q*�h�;���^�axF���ҙFn")�'� �V*5���Ud2 �6�5	p�ၞ��t�C�G�Ū���F@��'��OO�tk�����O1�]�q#������zH0
�3�
9@}���J-�:i⠍[�Z6&�Z(N�J���(�?wDM�&��T���Z>�J�Bt��?"4���U��%8�Q�+�}�l&o��Wd�����J>���w=r~�(�mV�ﭑ�:܄�Q�Sǲ����{A� �F�Yְ(���u�LԊ\�u}e�E��/�Θ�qZ� X�{���;)a&p�����W��ǹ��R3[3w�J�o9P:8:�K��m�J�������8~8'�>_���&��� �<���uơQ-�؝� ����~����|F��*�n��I�1�a]�H�4��p��b�6��֠T�D*J�B@c�Xn��]��Bp�)QC�g� n��>��8J���8�OŸNyb������?e�fb�m):2ԯ���w3Xd��|$eK��3B��F%X
�2M��[�_���(*w����L&��c�Xc������Wl'��2�g4����DwI��
��<�M.ҁ�nO�����Q������8ո��D0����B�e��/��wY�~eb2�V@s�LQ范��$c�U�eZ��I��o�@R^ƾ4f�0#O��%�V@.0�y�\+�	�@���+���~���8��{"z(��d2�����j�E���}%�Q���Za ?�����S8���� �A/�HXj~��w�S�a�p�?@s兪�ɂ�� h,H�z�xsˇM�g1�H ��b*h�ԓ��+���$���甈�@�V��
XX���	��Լ�^�6�s�r���zS>ty�L{���+�\��-,d���br䏝��߄-3���6CN�(_)��FEg�״�z�PJ1��@S�"���h��0G���Xp���<u�i���&�nў. =E�v���eo�D��{-�$�+�H�0�`�s.�NBL��>�� ����C�(��&2W��j�C��~��8j�=�M�(�خ+���=��r�m�/�'�(�l��<��y9���0�k��=#��I6���9=��u �2���Q�{>��g����!�rj&�Ⱥ�/�J�]���ut�"�0l��!��*�°R�E���>A�S;��o�����潣�26Vp_< kӌ��T��Ǵ��C��T�)�%�����dI���Xkv���kő�!�Oiz��㣵!�aZ��t��`������<���}�7IJ
s�Ou������d�d5���!0s,�[)N�@�����#w6����R�g+E���������7�\
���@��g�zsMkR���Tp���i:�鲤$���ݷ�/���s���h˥��ѝ�f]W�� �gb&��V)2Jl�!�L"] ���^�;�f�\���O-�d�k0���h�����_��}��Usi3B�t�Y�A��Y.�����1�ol��(ņ�-�m�'M!��+���8�Mu�<e���g��^}!�;о�yU[]�	ַT����[�&C��	��Ңp�4@�G���(�{V��̔\�L�ƾ#�o�2�y�Q�g�s[�,:%�smþ@�m-���<Y�˸r'S�]3��w��Ze�^�Zq�p֑��썎�[���q{�t��7eA[���y��A�?$�:�9���J����eu0p��שa�y6�cĔa?Q�!�H�B��&��b�E�p�*������7Vc��/�f��$���Mo���9�O
�I��� n6��Oh�q�]�	;��8��N��y�2?��\����wIu|�9�TG�^��� ���X���a���\͞�^��h�s��1��SIXiC��	��t�)b�K�_��E���J�UP�x��+�^ }HM�����F&gÿ�㩒���WO	��\� \�5Fz\��"�E�� $A��K󥥔���9��5�ܧ���=�}뇗�v�װN��C�1�)(�d�6��N�%=��&���L�����{~���։�#k�x=�²�m�?��:,f^���(�J�MA�ݳ�Bg�p6b��
a�`��%]��r⟉�:l����[&x�ʉ�E��:E�S��!Mk���c�(�ޞ�G��C����"�=	�&ig��&	��z+�1e��&�󁁿�"s�������|��Y��,X~]`��Q7��;���0�G2K�p�;��*Z�V	�0�k�2}���Ԇ��K��`O�;��J+qȑ��p~y��#H,�t�`�ԭ�;��.�׃�ņ�3����C�_��k�!Ѹ��݇�zNG��IM��PF�oW�K-1��Y�'<�{�^S�Y�x?�B�� �&��ҵ�^x�(� )�J�B���mm�1�B?��̕}�����|" 5p缣a��#��~)�-���%[��I�/�W���^TY�ޟN9����q�id�g}��ߤ�D[fG��lV
_�����j��iG����5��lT�Q����ť'�v�I��3������N�0�ex��*�a���x�0��j��2$DKi �r���+8S^.��}/{���9��.�	���[�(�2�(�L�+'��$>�I�g�"Y̦zH�7Ux�
m��ȟ���'q��� >�-�)�$i<֯��}׀2&�bw��$6��p��VF���� k����EO%�c!n�>u"���|N�a�Ҍ��/W琢��W~'��Zf��5(��L�,-�b��bl�2[��O4Q_�m�Πx��������n����-�j�lP!�Uͷ�$<��/��U�mA	7��u-lrS5��%���k:�	=��~�o�Z���-����iP-�`�|���������y;���:`�_��� d*?.%���EX�ϡؐ#D�C$�����[S;�z#��}|����]�ⴁWZ+��CYb1�n�6���9pA�2��Z-� �άK9�y o�Qk7���������y\��*�i����5������y}�m�s�<OE�;�)����hv�����{�D�l�N�I��1�a�#&�*5�X@��S F���|RD���P�ч<�O�B,5{�r!�O$XB�[��/�ЉY!��,�K?Ӊ<��$��)� 8�+�}=,�.|�cȲ��G�}�s�H� �!@y���ctz�'O�,�k�ť4M"3���{��"���m����O{~�'�E�c����d�����c�P�j�HR���U����/���O<��k�fl�ٰ�j�2_ "���6�Yej�+D����N��;T��!�(.O')J6h���=����\*�r��'ݐ���T(�O�61���E�%�C���O�l�{����#h<x����.�O�ZK�H�����̜��ڲy#6I��v; ��P��������|pNr[�$[������S�hx0�=\�^�/�rp�v����ϑ٦U6Ї;�%y\���`���I�Eu�7f�,P�R��'
<�){8.L?ʨe �1�ح;9��&�x1��3��Rœ�B:9�"�P��ϴWc������͏�����N8���IT)z���Jx�$N{�G���jܾ��~�� U�p�@�qk�ŉ��د���)�N�ӿ�ɬ��(��G{/=�*��ơ5���KrRm�%O(rfs��u�%o�oL���y-ӧ��O��8w�"<�`	^���L"1j��Ŧe^,I��Dy�X.] F�P�����u�K?�ޞ>B�������	��Y�d��3��1;ޑ��4,�����S[��@�y��O����Q��L:gs�5��{ϐ��x�����Gc+��BEv�j_�%Ù8i:���sBK�!|z/xٔ���F>�U�f�r\ Eǌ���_^1��n4�ΐtqu�y�3��h����wԶ�=n���a\t�[���'/I/�W���E!�6CvB���s�>���8T�@�#L\_�(_�H�B+_sa�mK:
����j��H��E����(r��.H<�fB�A����5qx�K��d�ev߳B��W_��+%�EH�v�v�̆���>�����:�����*�V���Q#��>ɦ�-á��A��'0���cy���I]��w*��Ⱥ�
�l^,3��d��h_=xT�`�8rk.|/eM�P֟��yQ�>��"�&���G�x�-h�ea�.s�h�J���0�p��9��Ъ,0O�}�-9�F|-�:�xr)�Sqv؍���(r�HK�x�Vr�ѥ��&��OV�F�b�Vz�\~�f��c2K��|)�[]8������cE�|r�5���3�ڢ�*��=!�U��UQ�^bQ���Q�����<w")�Qq"_9�%�8�_V	ѷ������ �9�h�m�A�T�Ⱦ$n$��-�d|j0�KBAMaFd��{hQ�UÙ�����l՜�3��2s��k�"��>�}�A�a�/�Q�Y@�D�a�.���Ғ���@���5O��չ��v
C�^���#{UƁ��.�j������6��H~ͪ<�#�]Y}T�b�変�>y
<�}�J(�/㢧�Uh�g� D[ui�\�,xt�����ʂl�tϾ��Rl����(b,� "�^��yul�"۟Tc�.�9�*|�͑�msJ���y�]�EF�GD�g�2�L*����29��v��[ٽff������@`�&#��#�mT�G�
g9��0<�h+�<iN���j�j��I��#��gL*�K�g]���MO�s}�`����4�y\��G�|:�T�ˎ!�`u�E�iB���ub�A;	%,u�س�^)o���é���#K�.�<��0��.N-	�'35�|-)��ւ&t6W���ϠT8�Cd1*_dg�5��^��K8S�:z�T���q�����R�8� �����bd�$:�X��F����L���%7�S��K2mt3�i5ߥ���� ψ��ʑܶ��D/5�0F�wT�l�J_���B{D%������:�,~ͳ
��R?��)8�r����h4�z��$�8�L��j�Q�-��G�u �w ���{��4�����i+LH��\3�*�a�&˾�0�v�	c�
薒	懩���AZ4l��F�e�(@�7c�5�����+�J�5�a�����\)~��Ԇ�� ��>/K$�mY��
-���D�.I�ȡ^�j��]s�f��xa�Ң~fCH��1�m����U������`�k��˃@G	:�6�i+�K���ށ7A.���7.8h�.����� ��`6��O��/R2���ʸ"1
�����]�O�Xt{bUZ�����9�Vh��S6U��?�$�|%*Ս�K�z͒��|���1i�R�YmD��k6��B|���.�I.�\A����̔Ҋ���U�� �3o�{6�;�O�����W�X'���ކ.f���*N��./�%T�Ղw� � �����b�ˉ�SjcMH��h���@�2�Й�m��� ��\� �#�+E����^���� �l	�Q� E���Ϭ�r�k&d]�S_9��Ť�o%����Ol��#�����5@���md5��+�B ���N�Q~Y�{����V�����'��c�O�$��������1O��7��HAIc��T�S?��5��>^`Ha���7�ɦl6L���:T{8!,�	�ߐe����~�0�����2y��w�:(�^2�}[(p�&"�"6D!�t�(��p��S{�*Y�Y�R�EW��VS��Z�A�@^8$��V��Շ��e ��7��/N� 3N5�m�M����1���d��I5( r����g�-H�ϗ��������1W]�N���X�N���V�C:�:RFbz~]t��	�>	�����9Q��}�cz���2�󪬦AUX�]6����R��L]κSrB�����<~��R�����ޑ�pRc�8��A�Ze��KA�_��99G���	�Yy�g|wK�/��g�l�y�����9�|#��D��*�h��7&,BMR������ǾqɧdT�{�w*�%�IK�V�nf�Y� v��Bݔ]��Gh3L~ܟ�wk:�
a�׍��
_��sY��Xľ(����y�-ɮ�k�����.�BHG���xNzةt�:�� ��Kց��0��ì��c��*���}3"��me��ȵ;��B��I�Z��.[�]0d_�V�W!;"m�e����AFn,o�a�������8�m0��>(m�+k d��u|���ȝh!ݺ!jT�S�b\�����hX��tb�S�2��t�IE�~?��J�gg�'L��ᛮ�4��&{wTM]�҆1�p1"TJ���������v�Ӄ5�V����>Нn��*�RڶcX�)^Z��� ��ѫ����p��/���?�J�OKmE�	���&���22�5�vs�z�(��7��\����]��ﻄ}���{E���^^;�h�J��E?�yީ�/3`G���hk�U߽�5�{v	���WL�QB;��>�����@��?r�CBVJm��%}\�B9�>ם��Z˹�(xܐ�ī�qt|�T
�-���9JSK�x�0Wb��Q0	��N�Pi���j��4y�-���T2�<��XH�T�@�H*?���l<Kkj�6<����.���CQS_��Z�jg���:T7W� [5x�^�x=�#�d�f���\��t�,�����w䛏"���_�`��\�q_U^�nz����aDo4�a�X��ࣼ`8*e+ƾ&���Ψ�p�}���Z|�z,��2���6*\	���B�qqP/��`4@��ܮ���,S9�xŃ��!4Ҕ�e1#����3�Ȭ�l:|�2x���q�^��T"'�a�_��G�rJ��GA!	g���B���䫇�&,2:kPÛ�+����%h���
�%H�f�U�-��f�h�[�
�<^���a�; �'V�g�4RZ�k��)��2*%�m�;G���+[�a'�u�� qF3c!��nk�"��Ƞ�<�1��i�f��H�KY�.Ӥy[�'������./oN�#%����ъ����=����(޷��=R5������r4y�V.'K����Kx	�/��zǗŴ:y|���I��'���o���}oz�� cu��/-�'��n��W�4�}93���5jT����d�@<�Wp��%���i*����z\��t�"�t`��֞������$�Pؔ�Hi���q��>~��`�R��-x�70sZp���̰	i+��;�-ߑ�\�>#�Ͽm�,��HU��5W����;��M?F�_q��V$-�J�v3{Md��ղ����%�n��������OB*50Z���~L>6��|��i�e���$U����XC�1a��}{c1�/�9��1�KmP��i��a�w�f�F��O?��v�f"1%����a6ſV� �N!�a�bͶd&#V���?MGJ�_v3��t3���Xyv�mj���� ��1��F�� ߜY)���9���:~�\�ĸr�F��\�E���y��@R���v"Q�$?Xo�C<E�*A�x;�]
��-7m�U҄�}��i�Q:��f���e�r>Ǆ�G����a���9\�N��Wmp���5��B�$fF��bl�칒�~���)Ȫ�I�>�͠�O�@��c!ʬ��DOM��B����[�O��`�}Z�G�]g=5� ��~�@��V�(�}ޥX���e��_ɭ���T��{O+��	�g�uBJE��4�YG�ţ�d���xVl�i���$��"�K�C�5��%x�F�"L��@�R#�dIj��I(V��X"y��[��b��PR�a�
�X:�7>Pc��T
����m�m��&,	/���z�M��5E�as���|����x��<>#)زqD`�kU�I�rV���?x�r��CSP\}�$���-�L�$�������1X1"}���70ZW>H� ��X�t�M��� 7�x ��>ㅶ�|�M�U�3�e�#�rN'����G`����+,�f"�V`j>��󓴀`�N_ԄB�[i?!�j��dk��F��%[�L���;�a'oD�r��~���G��R��4�|v6����i��+��u�X��Ư�@P��c��B*@W�� ��xr�r~E��>��͢F>����eH^�e�=���<���#<�r���u��=Ey�_��D���Y��zB��k�����R�wfo�!%Wc?�Q�P�6��-S�1i^�Z{_v5�3���=�j�qo�����3�q!R20�4&.����Au�3�[p9�5�xV���Na��:�fa�E�[��6r�Ld1�j=�K�z��ݟ�ˆR��	<ǌh��ɗ��wT�?��E��Q�l���ȒS	�b�p�ؑ�KM��G���꓇%}3T�s;��"��
[;���$�8��o��y���Ŏ�7���Q����������(���j��6���-�Ya��)w�KbԱ���d	;�ƧB2V���eQ����_0��g���S�PdE��P'��]�a����-��T_7����Q'v����5[�	�cD��ŀ���USN1�#�}SrLM�D��U�{U��L�/k��i4��~�L2�+b�U�9�����.3��¨�/�6er1�œOp��֊R5��<����wY�)1��ꃃZ����%/M�p�]����: �4�,46�zU�N��٣�I���i
��&����͂������]XC����Fm��{�����J�%/쪣F���K��i�Rhz��E��S���z�F_^��B]�n����K&�۔�]B���m*A`�it�1�e�DG<g�󭜻��?�f�Su��
U�6��� J��Wt)�H��u�)7�52�IV�1Io��C#j{R�y,��y<��nt�[L)Q1�Ay��_�e#��P��f�Dp�ʨ�.t�,�H��*�m�Ţ�3�Mr[b0a���ڴ��cK��R�z��S.�6n~�T��^�A�à�+Kc$=�E�;���!�ۢ6YڗSă��`�D[�� �A�wkh�%���D��.bz ��:���u�����F���~UK\�R���?��n����'��c�^�a� TC1����c��Y� ޽��EI�nY: �uU�SA�Y):��6@n��v��E����� ��בnN���>��%"���2+�\���>�f��1�	��\�nN�k��C��My���l�^�1� F�v_��JO��N�Qɪ�/��0��:�e���OڂD���qX7:� 0]W����$����ã�YA3�[�{F}�����]_ǉb�6k�v�6��DLF�ߠIb�<�P<�=P��͘r��X��\�T�ޘ\C�u�EˆWF�Yxq�2/�DT81-џ�w�X�3����p��={�"���V��ח���%��^��v����NO�V3c��$=6���D�x�-	QDU�n��`{���@���\�������+��źN�1d���?��wSz��G>>�f��p˧��!�@z�vI��1�ۑ� �����MW˶�ұ��c�H�A�џ~���1W�k���&wՙ���Jw�3���K����ʐ���U�/��/�Jw���j� ͛U[�������YU]Y>[2���3�N&�:_��m�ЁG�����a/Ge�B�l����I�`8����6�"�aP�N��#��i��\[��pHGc�U���m� �-�#e�_Ewe#�x�mD�jl'd=PB`��pX#E��y`�7b,�t1�<m��v�)o��[]L���p#ö8���6-�@re^�~��(������UmgёaYpL���Ʊ�fg��LB� Bl�3pn�^>�'r$�r���1?�顖܏��`�l�5/SL�x�IM�@L]9|���$���޼���%h�uϤlR,�xt�jԐ����}b�Y͟�;�__�r��:�S����X�⃮��ý��-����v�b�;NyƯ%��c�[I�|N@�tp���a����B��S�����?��'C�
�J�Ȟq#3Q�IzK��U����SÔ�~��ʜ��	��S��h>$��x�ZOKj����g�~©:�t�&��ݟ�f�n�� ����Vs��@͏7*MHp���4��~�#jĬ�s�5i}PP,�CDZ��=~+��(���Q+�ז�g݋�!����%����h�mB���j�UZ�u�ZR�.�{맓g�uƆ����c��q�݉ʃQ$z�4��۔�h�����*X�Z�-k���\�l�`��@ޔ��!`�'�5�i�p鞕?���r����nj��t� ��^���쌅�*��90Ge{��r�%I��z5�������W^3�3�Ά�c�1$�l�h�qo�3\�Ϥ���"��é�8=:F��[���!��oĻ��rq�gk���GT���\NvQ�OfW�g�5����
�сU���V�V8�ns�g}��n;<$h���V���*
�Z؊��J��z�e	Bn�v�!F�`#M�����|�옰�K �K�5q�gf�Ȝ9�]E���r\H�_��*�i����1�0Gp[tNTDvXLd鹐�1b&~h�`��#�9�) �&���ƚ�؃�H����?��ا��)��Na��l=��m��,Pu���o�����!�htԟ���ـ.f�) Q�A���G�Z����_�x8�\�qƗ��>��.�e���?G��CUK!ͦ��	\W��V�{uӁ��+w	�մ?;���!�ɖ��{��ߡd9��F]O,&WQnΡ�P
e�>�?5��Mlհ�4��Z?�1�`��l��s\���h����g@�0E3�Ř�ǀ�5*�T9�Ư>����M���Wւ���	�)c�_��E����4��;��`}3gDG&�gR�����Hp)�m�4�82�7<�p�w�$鰧�X�-�x�4�K}���y�:�B �Bo۴�0]��06�M�X	�i_D�a{��M"�r.��w2����y�$�^���R��p
A�:����?IiEJ3o�)�K �H�]Qd�6O�C�w9hF�۲�����=��HP��%Q�5��yc�⋝��UH��V���졙m[��^�<�O���o�P������}��T$&�c�*u7R.S�/U�QD�[�����EAbX?K�a���|y���_(�Ӝ:.�׼�e���oC���U��@@w=b�����dT�-A ��|F}�p�+r��Q���{�b&�i��f� �U�K?��Rkv�Fлᐟu�I�ok��	�[�a3x_GZ�"u��_ʔUF���"�_�&k����I]���?�0l����<dl�� ��28���*��N��� p���@7HH�|�}A�4+�C�]J �RO�!�8/��9{b�O�(���^��ӯ� �9m��; F����� ��0�ZH����I��`�����+����y^Ɖ�u\�y�N)}��6T������
�Y��H-�Ŀ�k�Y�/w�7�#�ʐ��ao���N��9��%���� �0&�`g��F��C�9�� �Ӕ�܎���"f�R�z�Ca��#Q�����E��Gb�.��L5~[��Lǎ3F�L�§�����J�<����{ݩx�T����լ/,Sa%Wm�sz�����U�;6mE�4j"IN! >��n���;uo�J�l�<�o�s����j�$�_��ȋ�C����KS��Fc�?�{Su�ou�&�����oK�M�;C���y�{��iܮ�G%�a$A�/]�E?��.(�2�s�|uxm��i��ً{{z�ISe{oy�1��*�*�Ӧ��|db�?����\�{����3�MP�Vm���Le��y!�69ѬS��w����&�������{��݂٢���x$��_�
�Lɫ�&��4�U�V��MetYV�m.�pE��)E�h���b�V��e_6�@IhI�K;.��͇��O����m��	r��B�V�=�A���,��juk��s�\p,���&`�b��&,�j!a�)�Ic�o�F�1N0���ؙ��l�I]:(u`x������Cf��*6�����#��R$i+��_HϥQ�`�R���6dP]�6]v�x�!r�kO���UN�Flֵ"�T�����iF���IƗ�1���9���f����Hݳ��1֏hw�`g�AA�*Lb4tn�8T����A���n�� o�E��a��m0��c���-B�v�;l&n\&h��y�ٵ���D�hcq����f�m��6*!M���x��R�I^�����D�G(��B�_yg1����b397�d�{�^�*�h��ǀBv��D '?�u�OF�Wi�!Au�4����\�GZ�?k@?�-]��u�X)���o)cE`O��� 
þ����G-͑��>/`�b�5?�7ۣ�4XZ�����ܧ-@#�X��t�8�k���Ҽ����00mbM�_����Ajs�g�#���il�����(�p^��}��n$���9��D�b�_����\\"��G���C�R��|$�Pc���▲>�� 8�3GzFqSz`��x��W_5���@uU�������ݸ�E.�����^��v��&�.�i��1�'��~���ZM� ��i�������Si�q��l�mӔ\jk�	��5u,��Ӣ}��Lb�t.�6$� lO�"�:+o^�1�Q�E.�4����� �}�UP(4�`��)����}��� ߦM3�š����Ǻ"�Ot�B�H���yj�3S׳����7�{�q��kİq���ί�6pMD�7�y���l�&���E��v�wu,�1H�#	�5�冺��Y�/a��9x��U�����|}��\������	ψ��L4��Ο˯��]w\��~�'��* ���+8�t��I$Q�g���4�w ����|'��Qb.�/g�n9vS/7�����BX�d�)����Q�X3}��`�7
��Yo-��^�K�#��$|]���M���j@F��G�"&Iok����E���P�i�ePM:7��:����q��,�d�ρM�&���D,�~)�ޭl�R�I.��M�Jw� �ඣ�g����3����" ,��p'�z�S���y��C~b��R=υc[�E^(	{BD�ekH��jP;��������8�N���ys��n�I�g�`Z�����J �CЩ����_�`4Wh������8z����#QGz�9��V�C>��Wq?�]��V$���}���a�^���;=�Y��PP���ڌ���i�ӂ0��>0����E�=��qah�i���?��f�"��K8�z�0���!�
��f~�7��@�N��kƄ�p�C�C|�ɸ�y����0��YE��v��R>��W9�H�io�WǸWd��Ƒ�<F�!:�����~�� ^���ȓ��B������j�^ٺ�f-�ї<���@䌒�T-A>�!��1��*@�Q��?��������\��u(����h�t��p}Od	 5�L�z��Cr����	��k�(��I��D�xS&����}�q�x�_����+��3��}����h�\%�p��r�����1�bq���f"{[���� �ؔ��sb�_O�(�͠T��?	�Ǻ]ƣ���	�Ӄ�4Մ895#������Y�.1���'�5�ѵ���g���6���'��tU�j�ۖ5g���N�)�o!#��ɘc�J��㘜<if�C��e��Db�ws�_�r�D庀������๦��I+�ң�:(�3p�� ?�bk��G��e�0s����L�ݟ�����-����a֜{��u�`�xB�W�kV�CȰ�m��Fm���'�� �!OGK>���oWFD�F�V${�>��&}�g�pt�L�8.L��l�UA�?E���I�t;���v���P_`����M~{�Z�t�q�$"��-�A��C�lsR����K	�ca�v�qd�L�Ko��<9�E`�	ǵ��I=X{�C�����^�'�C��S�J�WA�F����\4�k��o���)��(�3@���({6irݝףW�l����⮑�RB�>@�O����B�Ԝ��r�l�v���_z�{�t��6	��[B�mF�+=����.�����1��f�-(��Vy�YWQ�y��*���~VxFXg��p���X�%��봭!b��=�Ab���^��_W�Ep���#��&w�O&�]���@��z+˜��$-�0M����¯�T]�uN�5�����;�e��k�@� ܔ�z��e����Da.��Xp����&�X�A�P��F��Ff��?S踠zh[�b5�J� �=�b L�?U��i9��#����ږ�m*t�J5�@�q�ɥs�T����]s����b͘��[׽�E�&[oh�xc=y���0I�+5�S�@���n�jx�,�¾��������m/�Q����]qx���`)�����9�$��Npv�v�;S(��X��5���ǐ�����v|��޿���W��JE��*\E���1�$�X`��A�8��M%�7|~zo�]�u�h�����i�(�F9���{�$�z�:v*�(巺lp`��tD
!Aa�$��خ*�)Ș���Ƽ��gH��Ӭ�{��Q�8�c݁��m�ňg�b��g��Y��YNx��6%���~ײ�u7i�M�?�ks�p.6�5rI�����0����m���>��:1�)���}=g Cg9�w�����Q&Ɓ#��hh 5�C3.ƪ��˔��M���O�ߗy��s�Sp����t3�m
Z�8`�!3��0�n!��}�����<u-���ș9���[Cr���L�/2VA���� wt/^�m�E!���JC'A�ٝ�z�q=�P~L��?��,��>��m,���O���;d[�b�d�vR��E�Q�%q���p�*�����ɜ�u��w�� ������jX�^�j���~�r�w�k8RqB�jA$�X�Wp_�1���aZu{�6b�M���>1UGC���C�脍�12�*���vi�g~���ehƕ��UTD�5^e���8���2�ڎ�o�PR���#�3l����k�P>��k�֮k���O#�bs���܁޵��.4��4��-�2y!*��A���fPX��ҏ�xBi���LElU��P�(�p�>�:.��A��Fc4x�E]~(VuzOKi�/��@qf������C�@2!;j�{�k�>�h�	X_c��4�.�$�[����A��V_"6�.�Ѻ)Z��y7Pd�2�!���5j"�"��1�nqgrf�����y�Ff��gp[������b��1+��;6aM�������?����Xq}�����8�6�(r�M�m���W~��N,��%��$��-��Cxe�8�d�=�.S� ٸ��t' ���)�yz��s_��r]p�`�\d5,=Ft`Ϛ��r���%��sagy%;_����YG�IE������~p�2S�L䳭��R^��_�F�W?#/	7J��]�R%��¼#�I�I�8p�ƽ9��`#�֟���8�h�(�����u�]=�
3�EF��=Mt&��77��������)m/��:��i���2��H�s�h�C��LN%^�.I����rn�_� Ô�Ϯ����+d��qE��PH�C�Ͻj�<zK�%�.���]͞�O� ==vڜyR�
�@1}�T���B�BKФ�D[��Cw��9^r,�I�嶛xv�(��\N�ގ����5�)��E^Und[,��(��G/q������Rwp�l��^]�듥�E��1�iK��H�I�2�Ju�i�_l,�� t�5kʂ�{���S@���`��,AD��<O[<:?$�WtB��kභ7Z.�LXeJ�W�A3�aNC��$`Z���%�**㠰�Fp��wۦ�М{�T2�}9} r1�r�EvQ��վA�=z{�L��?BqPy+{��O����ѺU'4IEHF�Od�ٗ��X?e0�����zsK�{J���0dG~��0��|774~3o$�ڕ+X�j�+�^<0غ	U�:0��ՎGa���7E��]��q��o�G�d�y��ߐ��"��T5�JM��)�ͧ�h�����}����ݽ%��}��ܳZ�#3gm.VT��;^�v�}��NRy�m��o�5��c��>���v]�H�!cG
�H~T��Ӂ�+Q�J.��\H�i�>�i�bL����������,�T5���)�yO�?�����Xr������ϐרw�c�.�Ut�?�
O���l?`U������~(+�p	Ju�@����R~#QG���M�g�
F,�Dp��$X�j�.UBUc�:٢����cL�����x�>n'+�j�^��cfz3��魣���<-�3�	E�"���Y}���Ao;�fV�����2MPפ�h�nPs�K:�O�e���H�����*���Rm��hn��˛�	0��3�T4׈�U�laJ>o��~�۷sٞ|@ gTl.$	t��=��7�	�Z7!8��>��	�~�Dۆ��h��+n!���ZxC?��C �[
m�'��`Fڕ@��B�t}�2��/��;�K%�f2��0�,�ӯ~$�{bu����iȲW�b��������c�S��>CR
ke�*Αѩ)��6����1�x��A���z|dv�-PLZ`��4�ઌPo�5���'~+�Z��S2ߴup- ��2db��z�Fޤm��e Q�m��F����:�ã���KXY�'��^:�
� >�X���I�k6L��y�E�:�O�7���|:��U��3�Dہ��ǔp��<f��$�Az�e��ki)�O�[��-�{8$��ҍ��	�О��yn!�~bK��2���V�H�}׍gs�c��[So՘�H�B��i�RMcH=_^��T5���L]v`e��n3��H������d�Tu/�+~r�1_�=Q��S,��'2M�&�]+Q�@�髁�1����&n��F�w4nɞ�,�CW���F� rmE� �.�Cr����#���|u��%��ȍ��S�-�]]?�>�Y��<^v`o�;P<6���2|�?� )�ϐ0ɕ��i��j�N�z�=�~�q����"1jh��3}r)Mȴ���)��� �e���^���Iv�1�:/��^1��S�VS{�9��d9������T�ೊ:� ���a5rj�I���W�O&6 ����b�����u�k <*�L`��^�Qc��Ա�e�m����v�س��k�/�(�*[eWPBWP� r��Ʊ�i�����S+c`Ϣ�u��.7���V{���VU���^D����U����0����񌟖��Ƭ0P^���OԲ���WX�ؔw������Kz��6��0Ǹ<�	�:�^f���E��o�����8��6r��j2�gkP�j��V��.A���j ����=9�Ԅ���2��F��$g��)���;a}�_�4�y5l��%�i\��"Z����^��I��jB����"*��[J;�� �j�:����)1ӳ#j%{�u�[DJc|�J]�.R sjof� |�"K�y��f4N�,:ò�+=!&�ma�P]<٪;��':�1*�AC&�H�q�	�<-�]��� ES���$1�"
GT��!�Cy�b�(�dޓ���;i��	 X��h�$�F�*��B�c9	y������FkA9,ZvM�gil.)z�,<|�p@&����|]M����:���Q�l����m%�}W��R��9����#�)a�!-��*G�}#���1���)��ɭGʱ�1u|Z2
n(��>����OP>a^��U�c�h���8��\�����)�2�Ń�ӱtK"�a����X����"}�qS�,�F��]xon�EXa���7�74�N�uA��3�~,�(+vܬ��e���܊D��rb���96�Y*U�v
|���AĻ��NX����-��uǘ/�Y��&� ���A�'�����Y������v�A�]���YX��	��-��mƚ?qħJX���}��I߾E��w�E=S��6L�{��r�;��iI��}��	�{�U�'-AcG�s�ΰ�ӷ�A�{V)$7�l���
&�$�H�5�h�X讆y�o-�rc�9c^԰�'�g�1\�87p�ټq�� �,�?G�?�&i.�c}�~xϴ0|�.h��#����){�>G47�G$k���h={;ȹKQ��"�'!{Z4n�����F���j����������0D�'�рُs�[��̓��Z8;��}J𖋁�T���<6�V��l�)���ګ�A�;R�T��#-ਵ�*Xt�6K�[Ms�_���l�y8���H���$s_���?���f𺤌^�&���P����<E��v#�)��i�6`��~g���%)Rޢ��l�~i4�1�|�� j�py�n�!����U�>m[S����}������G9)���0��6�CJA�U�B��=w��OYu�'��&?#�h�
���M�eM:�(jՐ
�=���uܒ��ѮT�x�<��ޘ����0P=��x�-L�F\#m�9.d��<t�<��%����h��q:��*_�kc�Q�0S<��@�i��@h�V���-��:,r:�{��/�������5���W�^ҭ����$�9�Z@�+ű�6e�յ�����79���#ל%R��^����L�sc<�=_��ՕB\�u$���W�>׾y���0k�G)��f�J�Qȁ�����Vm�����Q�Zn��`�Yв����7sp�B�MVt����e�æ���ض_��97p"vrA�*��и<���D��I�W�e���O�9i��*��];%'����IbfW"��N�����d��o��we(ͽ�&d�%Ԏjc�������>+�1�ߙ�@JY�p�:h�F!-�������3��4;�K�u"���@��1k�ژ�R���؟�B�e5�4�BjO�o��}4#�*	)���'��e�_D�j�hsW%��<}]1Q̮ �� %%rJ9�"щC#�����"Wi>�L(@�����XB�{�c#K�d��DvuAc$΢�-�ً�(b�������3h�gqӍ#>4��:ے'cFɱ�_9gn���K:m�E!9V��/@��z'�ʃe��ŀ2V�(����'�s1P c�h�ڱ� �d��<䱣���������4�mj���ܓ��y�%�7ժ�C����7l\��^��%�����e7II�����RE�_���[�n=����}��Y���qQ�����ZCs�m�HJ�k�[�{a����b�ͬ�B�S#�zZ vA	���܈BFl���~��zk�����z-�b�Gz��9�:��JX�"�-OG\����&zB铗
��E�,�B�!o�������voC��p��rV��:[�E,��6����k����j��[Po���������(�5/k���CrbH�f`�,�o�EJ�����m$J����/�1d1� ��� ����)�}�{��CN�!M����MQ� ��4q p9"�X�gg��9�.wK��Se>:P=��EP~B�����{�ؑ6&-R*7}�唤>�L�s�t;��ё�H�_�b( =��{[h��²����2�N;�p���u�(˜IA�x0A$Q�Ҽ�i���_m,��ɺ��예6��BBID�L\گ�IŤ��k��"X�ҁ$31)������9����l	���y]5Y�TsJ��y_ך���"�ݠ�Y����aWÅkc�0�fm��~Ɓ�BgG�>%sт��!m��4�V5���m9.�3�ω�Q�k��=�J��h8����;��뙄5�E�D��Z�'x�<@�{X઻V ��Y�D�'�&�U����P#�|^	8^��Qx�4}����a��]����q�G����8��q��rQ>��Yp�7�aҬX��M��E�%��Y�0ѷ�w��;V� ��q:�n���4���4+�CE��+�y R�����5�*�?M�|�@�(�X�y�u���T�!t��X���/�����t�}:nd����"l�b%�:�L�hՋ<TD�'��=;��{�ݒ�8�%"�rNlI���=�1b���v�9��G��R���0Y
�Q�U
Hj?Z��=�qt0S��)ߺ9��^�K���#��\蟐��2F�b��������܊[۱������6��ҳ5�FD�I�2�pazvz���7�~�脵q&����{  ���x�7[�1
{�r�	?ʜ~g���	U��$7���[z-'�O�X8D
^��Q������͡��
K���E�!��d$� �<�Yt۩�'�)8r��뼅/��"x��U��D�g�:t�L����!R��	�ܱZ�pc������;��:C����XRR�C~X�T9,IX�V	3*;u� sҿz��!�i@e�|Fhu���q�4�o��b���	{l��=��O���dӐ'���b�+�q��_����+�hp�Ҫ2����+7F�A��{21��3�`G(aB$=iYV��R���V��q�`a�cV�`��J?�_�r�� elm�W7��m���eU���s�o�)�=�8�~�VO�U�
��(�	tt�����"e?��ns�ӱ�/շ�v^��/�.n�$�N�$�d�SP�z.�vrF�����wR+Wsɡ|��g��.�h�U4�ϫ�Q:��}�)Ro�7��\�sM�S~��_tr��|�f�QZ�J�ᘸ`�'��<j[R��H%�AG��	.ؓ ��I݇�_:M�D9<�hw},������P�bRG��8w0KF:-ɀR猽��b�~�� �B�`��,)]Bh�:>h�n�#P�l�9�pJ��A������T)
I�`!���M)�Yf4�{09͞�L��_�Oۇ'���7��d��a`��0W���k�J^_G6D�]���j���V����D�Įc��k��(����[�b�X4'Jp�L�GD�_FՌ�Y����۵�-Ƭv:��]�H����gشف�kּ�B�D��/��O���⾣N�Ր��4�����		��^m�N��9m��f~����Ƹ˅��3������ӸiX���N�)fr�vI"��y~?����Z�l棵gp������/4Ԭ��|�U��աc��~M6M�. B��KL�P1ݦ��?��h�Sy[/!�Ǥ	�$��m�U؄�o�w�5L�51�B��x5���{�w�ی1�s92��'�{����N�l��+�R�bm���r�C`�y7�"���޺�i�j*Sz�3v��ֵ'��4n
��v�K�JQ��bp������
D��VycE�y�SHB�y/fU�һ	mz�`��HJN���v�!"��`�[6�Gh��n��1M�� ��t`���\ff�,���Spg�8?���ǌ<��?sXj��=K*��[��0��&��X��f/(˾���¯K[K�7����X�?�0�۽��E�!X 썩md��_�՗�1�G���56�@��47��Rt����$ޢh���{<۝�����C:&��ID�/X6��W��6L�z5+��{��o���e�F�fͿ^rS�Q�V�����Q�	���d%GR�j��S���}��H��w�����,xo�F��$Ƽ�No9��*�ǝ[� �i)L摙��Ѽ{M�as�������.F*������8�I�E�Xa��� ��$:��ִ�).��@D��lH��(}/"� �Q����DE!��8&`F	�����Z�ĕ�߾�V�t)B���Ȳ�����Z��E�=#f����[�~.T�Q\�]�4A�=_�,!ǽ���pM~	�|=�8�^��mO����5��Pi�v�%�`n5��0@/:6CRE��%�^g��$3.�̗k������;F#������r��B2&��!�fE�pDm��;�vP�_�W�����i��Qc���2��ʜ]��eH��O6��{�k�ɥC�[+�1��d�����mK���UMuD�p����4}��u��v��B�Ca��'uɏ}�:�z)�
�Iо��5��
��@��=A�$�o�lb��\0���YEo�]OQ�	qSw߫���nY+��(�9�iF��y��k�R$��}��݌��$����݃����Q�0�v"c��;�7_�9��.�ژRrF�e� }G�]���l��xJ �&�qP=������Y�+NdЋ'<d�K�#��]��5��`�2I�|���v��}���|����U�7�+s�!9�}�2�h;�<ʘv�J��]x�|P���t����z��gҥ�}��A�[p�$��]˳1-��˛���}��$`!(�v�Vh>�8�c��#��:'�ی ���m�U96=>z5���V�x��|��G"����/�iO�gVuXg���g����������n�������A��!%�O��K�N���WM}�X��t/%ga�~}�%��Ps�����Y��x��4-E7�T�Ic�R�M�Z���?��5�ݫ����/����FC�J6tC()p}c%jyd��O���E�4,���)�QoMG�����qQTy�%�M\�M>d�ʢ����$fE?Hh}Ä���4�}z��Ӎ���\*m�o'on�a�R����,���'�E�uw������$Կ�|��:\8ؘΤ= ��GBg���㰪3�c3fz~�z�x�t�U��D��@�6� ���!�xqpa��8P󳨹R5�kÆ��;o��+Iٶ	�����m��hr�F��X��}Np���xh�(�9�I���󼽘E9f>uM3E�0����v,0�����PQ/C�;V6��l"�3�%ēy�W#���	!�eM4s�_�R
+I<���#��E����Mô�ִ���%�#_G:��]�<z5��^d]Xg˵m�Pۑ��|��j�w��L�q�źI].�"!��u}��.��9����c ��T��_��rI��Ί�'�T��.�M��hwƛ|¡��T�e����A�{R�&c3��Iu�.�ӑ�l���w��� ^�k���
52 ��B ;b���T~!�y{42�W�Fzjy�Y�C
�����${�L`4�g��>�+��6;�lE ���J-U�K�X9�R��Rb9���d���Y/܂0N�q�C��9�X>���]�IL|����Ju�S������H�يd��W�Ӕ�W=`�}rGr@�bS��/�8dU����a��d�Y!�9�5�5�V�><`g��b!���Q���剫�(�Ή��*���P�-SO��*3�ͺsy��&{)[��&ɀ��B*j�G:�M��M#}����j��f振�o��eP{v�d��{$9�/ɢ<)2�K��H�,h%,9bD�#����? �*iS>����Y��:�'G3��*[�.8f�b�i+w�{�5��.���L���'�nIOE]��1&O�>t7I6�J�̖���|���#̀�����>G]��?V�X�-��		��(���Po�9��n�p@�-��tۅ�Լ�ǒ|�F]?`�} Ak�Pk�\ܸ��SF�.������y�!���+E���*-�fO\Q�!�̬��F�{S�Q|�\.Yq���k�]�8W�rP�)��d����ߝ�|D¯�N�i�������psN�R�d{���E�~������Np�8�#���G��̹��\�Y���j��i�j.i0��>�=��%�n/���k�o_UN��)4��K~�$���i;θ̞�w��Zc����?�������1y��Dp9\E�*
���4��<�4��KZ��[�`��9�傂�.���J��t�%���U�ɖ�~9�Ŕ�eN��Mn�}��D#�l��$r�{�+�x�VG�w�Bh:���� l�`�}�XX�d	���Mr.��J��f��8t���q���l�/b��5@_�G�.XS��u��&�U}�,�qа|�م/3a�~��C�_��a���R�-������t��Ll���3	��Å�𪔽C:V%�~o��A��pV��~O#8��.Y��{>�r4�o@?��{dc��'|����3 ���fhk���%��J�p�qn��&u�Y�O��� OW���)��ID�%Z�8=��(l��1��"�O؜�Z�T�o��U�-,2ۭ�j�g!��?���C:4Vr�^��N(���(�<�� ��%<�yFkV��.ٕ� �(��/�{
�Ւ����%g�zū�Xz���d��o��g�4��&w	rJ �E.m\�P�mc��$!�b�`I�O��9LԄ!�1��9�ť�i�����H�#�`��k1�y͚�wo֝��(a�HW]�l�I�#�ۆ�э��p��s���1#��Km��ڒ�t���(�Ցz�bb?�L�8s����2tu0����UB��l�	 ��� nt"���FNl�g�%]5o�o�V�P�0�ԎZR�.��92!�-s�gA1�f��b��	)���W��A�6 �5���?<��O��Z���9�Dǵ,k�u?]���R�~��3o�.;����0+B�ZrC�����`��%t�Sju�吹� �RH�g��Y6�F��0�
*Zx�ES�Ԑ�]ܢi��_N٭Z�̋D�p�x6��#�!۳w�g�#�6`u���A�b���d|,�R>_�w�~=�U�̈́�'��O}��ZmU��-�{��jb=����%Z(�?;�o�h�٫$��SI_!+�I)l�F)���kt�4C�]OOa��)j���=���ص��}�Umwa~H�C0�k�n�q�C�PI��$�l+��	���N(�U�W�}eAT����x�-��e��U%�����0�|�'��fH&B����7�S��_��.�h-?hvěA( �Q٢酵�3���o:�+��j����g��5��/������~>���[Z�&6޿�V��
��
�s �K&)1�f �ʅc��q둃3;�z�%rbz�vtfJ��y5W�Z����
�z��O���� ����Qy�A����J��t� Ty��px�R/��qЭ�^P�5�N,���Z�ِl����l�o
�" ��#��q%԰��̼,��'�"�EK��Ɨɂ2�%��ɍf7U#����ak��?��_!lzHOq$XIM�]Jx�x#�,x�?��g�Ȳà�d�:n��)D��'!�#d�~̓b����b+w#5���3�}w׶(��tu�?��QE9�VȬ5������"��
kU�a\W��+�� ��<\-jZ�\^r���A<���f�1כ��h��P�P����p5t-:�����i4�8�&�5]�f�<e���T����� ���\��#z5���B֫`�	Q��d�kE���k��X�0��+�ɷq��;-4��>��Y��
3���D:���1qb�ZD��P�$n�9��Ȣ���˘Ț�L�~o?.)����j]�8\��.{-^���r����X���b�n5�H�\K	DˏSY���2���\�Cdeuuw�ӆ�%+ ��m[��I?
�lfQ
I^,� ��� �l^�6j�u��>#�fv<�9]��j������.����$`��˽��e𐣛�#���$P����T8ߖB�9���!��BMu�7�1tXJ�0�$��m��K�$��[�S�^W�� �*2c�D��D�Z9�4dv���Jw�|�<;����O#6��ت[c��"M t=8|}jQMM�1Gc F���F�4�6̷��s2�F�-9��@�Lώ�ET���m$����j]&��V�-�ݤ��m�A*���EK��8mA����#��}�@{��z_����0㐹&��Pi��G���YTRg1����Cq�T_��(Z�����^��d$�_Z��s@�������҆��X-���awbV�n�2~+�u`-T	�t�w�G5���b����7u���h�Y�����E\�0M��x8z(�mt��@,}�4��Y�������|mP�fB�ex�Kkc�i�K6���Z���fY�dW��ؑ1�i.��9wZ�I9�TL��y�ֽ;5��)oz�l��\����j�Æ�\z+V��Y��%g�<��[:rl��\硄,��Z��Q�^����~���~��ZR�jo�a��gp�X�����s8���ғr��|'�_QvHv2�M�`��kYN)��5��@�qxd��0���q�D�T���<������+?�T���t�^T�|��o8�㖊�_]���Ñ��xI�Qa,���"y���S�+?85�a�9V	6CsP���	������1�Kz��Ԥ&N���A���$�7�������Jf�l�f��u�A3��'R�*��t(��m1Pa8��'����b<���%����kX�o�앂,��t��2Jحb�e{����>����i��5��,��|�w�T&���	��W�<��������D��ޙ��}�e7��^��o:n_s��G��X=	Ls��iN�P�R�9��i=�~�Y6 ��(�Q�s���f���W�Xb�iՠ��t4�0��ڿ��e�?O���y�
US���{�$�'�����J�}Ԍ}�^��?0IX-/GkJ1|X�+�n����V��Ê�ε,Vi������ ;pM�����k�@8�NX�(�#������ܳ/hhl����\[��[������k�ݍ�m�ҥ�Gy����ݵ��������0�A���`D�D��AZ�o������֐ؕh�����~����ң��s��u��a)g}b���t��c~QH�tm�c)���U�����T�U{B$lt���Y���y/�?��;'�~�k�d�a���G� �V�g�\��cq7Z��B[I�tFC�b�����z ���ӓ���o/a��M#�h�{�;ۿ�o��F?+���Zf�f�%��)�lI]S������WaY������F_x̯`��H��j��D���FK��×�
����S�e?X)�wddvw���g�7�%D�/�����E?	��ס�;-�.���]0^k���ׅ%��
� � �|cr�Kl��r�W��������[�1˺/�g��s�[̗Ĕ${���Z�A��t2�z�&����5,7ڱ�  �{-��c���Z�E��e3�u��jZ抉��������ˎE�Ǹ��_3���^�r�|r$'��V�7&N�i(��	r� ��8���c5�S�m���?�XMγ1,bz`V�?��'/���x��]J8b ���\}�A�[#t�
��� j:D��X@�t��5�	E��295�h�X�$l�.��ea*�8�a%����<����[Qx���,<
�@����`��2�a��R�}}_:��q�+0)7�|��ɕwE�?�/�'u�ƻ��e0JIۘџ��2,eB�/KЦ0����������D� �p�n	��Aɚe����]��8|��?�?U��B����#Y:PAMb�O����զ-�7Ғ�C
�O�Z��ig�A�{T�RZk�ǵ��xT��Qcâ�� ����o�ciK_xk=c��o���jT+��K����Zl�z8 `���@���������Ft�A��Jl@����j��C!�j5a�QM��ٸ�}������l�����~�vMp��WyVi�d�o�0>Tkg�h�r�� )��P!��͑����I�Vਾ�YSMy�E�O ?v��E���c��@�%�Y|�x�IB*�m{@d��Bd$l"
�vs�BZ��.1ƥ>�A��e�*�7���s.���ގ�P��e���m��]�P
da��+��Y��>��Lp�o�%ۂv	z7�&^&��]�[� mR�0qFWb�pw �>#e%��`�[����/3k@[&�>ξ9��k��~h���G��f��p�b7�5�.��]{�e���b�u2��:/?S����uu7m��s�s����Z�M2�M�f�#t��;kQd���~C&�h#����2'��q��|��t��fĉ������,ƣ�
�#�������@!���<+���!�3�/s�$4�@��: ��|��3�Z
�ēؔUmG{�>��w4�ԃ��?p��E=z��?)M#&%`�x��E.t����oh��I��:R�̬�K?ޜ�g���d߾�A���;�����ݒ6.]�
AX�O#�ub
�[<~�|�	��'��;|��f�mZ��ܩ�=1ƹ6~���<f���wƷ�ޭzS�7Z�V�� ��z�{���$���b���Q�z�U5�xP$���r��R�Ò���k��7%k��RK']��4�����g�(�m]�wD����t ȃ1@�}��c�b,|�j����bdI��n��R��&8�př���$i��T�]Ts ��N*|��}��P����ZJ)�a�}E����6�ŏ�E���	��K�P��� ���m�e)$ih�m��*�1�x�x��?��I�D8���\�]B݅���	�w�<��&�R����}���5u�	�׍���x�T|�8�^&��)��[�YRr$:ӊ����L�"���3�T���/�1�U/�S�,VG��iDi����me/���}��_�R˼w����V X��a�͢���9�q�1����&���sD�EfѤ��yؚ��xAyi�����MCYX/��j�$��Jf��W�@�}x�J0��M��֟�5V�`D�q��N�scz޵\���]�
�@\���ͭjǯ�A#�+j�������$�V��)��$-���gЧGnX�π����R�%���DA�n_��0�k��������?��D�)�\��[)�y���#㵳�Kl�YO
g��SҕlY)^2���iU��)��_Z�@w���+1Ǜ��}.PP��l7���ߕ����U�i�0�9�k�[eʫ��9(Y{�
_q�DA�YVd��J7�x�0��Q��	��߯�U�nr��3a�2Db����Lt�ބ[������0]q�3x�0�������V2ɤl����p��/��P��"7��5�&����ea����Ѵ�N;�����|^��M:���>^X� ��$�A"�:�F�\?���<���X7`%�U�D�9e�k!ڊ9z�Յ����M�_F�#㹚��C�=I�>����5��T��;�uet� ��XC�#��T\c��Ħ/U�=�G&fjȉ G�g��� 1)ge>��#�B��ɻ�Dn&�'<4%��S��O%O�YדFG����)N����Z_�Қ�əA�t�4�qڰE�����\n��]aV&]�M	ʼ��������?�[׮P3�x^፽%B6�){OR���^Q�}�G�ײſ� ��Ȅ���
Q@ q�ٕ`������HI�Gd�c���Ls�7}	C�����Pg	.�Xl�Fh �/6���������I�<�������K��}.yB�B�oc�y�����ѷd1�K|�.[�If!?ǃ���Η�	�ɸ��e��������ɔ *pֵ퐟�����'�8C��e���~i��)�͎����`�@7o��'&�_Ũߦ>�
8����R8Mv��~�N��w�E=��镀vu�)E��t���j�f�)�?Hs���Bg�BD�����
��]0n|*CA>�9��:�t�8Z^�@��I�(��L1�u$�Fe�e� ��k�-�6 ���h�hf�8�3?)�!�O�� ,D���e�E���l�yb��b��5��׮B�`�0/)\�А�%��i�kL�a���	�|ւy�n�B�>��n����G��W_����T"��[����[[t��*�O�b�dV��;��+I�Ϋ�U��c��Ǜ"H�=u��^1����l�tNz�N� ʈ��a���hˈ�a��)F-I�%���6(ڬ��vB6��bp�s��m!�,n$�����u�-�~Y<�ݰȴ~+� �Zv����YY�-��Bv�2 ���-);l�#����L#I��!��ew9�8�zv���[��:.��������L�݂���l�e�!�lt�t��!{@��	�(Kj�
���`��>�ꌂƒ����z�9Th�^C�����E����aA������Gr=ȹ����߷��P��6�Bw�K���+A���ǻ�t Ӓ�-�����{ʓ��B;�z}�������->M�y�H��R��p�t����{	�� ���hӶ��X�,k���#g�x;�&����>9(z3SˠrD��Η6O�/�J�9@�b�0k~����"��'�\5�SV(l}�����k>޾�['+�X����m��t&���&#
y������1㩍�e̬/IJ�:x+����J���I��!72Rs.L(g+X�K����tFM���w��$ �S�p�g�e��E�ݏ���{��/�ͷpv����V�J�$@��O�����>U�8C ���I��Z��-��/����X���ki�pߌ�3���P.+��;Tl28�ahU�V������+ՕjG5�F#ƣ[�i�p-7<�q?u���j?�F�wŴC��Wף���r�����;�̓���.���A<�����9�F-��(�p0��帒O�[� |��3��Uҍ��
.Gn�ZRI_+�u�&��7=p�b��.�g�3|	Y{02C���o��7�e�7�����cCߧ��[���,�@8͏�*Vg�k�=�Ťv�Y}\�g� ���eH��8��W}�S��|Q+�Cp� �� �_���貱���`�m�hG����9U��O�j�Ka������1
8yg�j%� ��:��@A�:ȊJ�9�� w7|�J�Hp�H�dD`G����l`�9;��
��
���-S2�ѷOZ!O�TןC`��v���:y��Gi�W�a�����y��N���1Y��8�M���o$�U�������J$?�|y��&�
Q�������I����c�i���b�����\���Ʌ���LJ�ǐUÝ���դ���RN��ƪ�2��m(**��@~����.'/����ֻ͜�)3���qje������#t��^�f3s!~ۼH���Ak-3��o�9���ۧ�1������_T��6��)[��g�5؞��W/��f� �rl�y2�v ����[�p�׀�'zt��"�c�.�Ʃ�M�Ks�@߸�n�Q�a1���%���oLmm"�3�j�e��q_�]>c�FGNG����u]��z�w56<���Ul��>!����v��u��$���z�e|���R?�ަ��=x�y�{/c�0��a�N:�F�i�J�W>]j���0�9k��b��C3���"5�m+<_�aoB4�L,)��hO��荜�%�5>1N}�w&� ~��	����oX�o�3R�y��5[��Z#g�5���x�[%��fևS酴yj/���9/w�� -r�y[k�EUY�-�-�\V#͎853��(+t��S�yug3�2����C��>�F:��q�#�XRZ�ǂ#�>~2J�8,��?�{ĝ�ܘc3����,���Rb�hVE��a�}g��4�y�6p	�+w��K�N�QW%j���� �S�=�n޹Pp�rv/L���]�Q���o؞�K��|q#N���'���*�b`{����tWA���W:��3�fU(����Ϧ,uak�NÏ%;Z�sI\����l26f�.����?5"�ha�0��M���|���{����B�i'�󋑁�Z_o�:�L�[jK��������.-I4U� d.i�_�3�J�Ʒ�<��t��ߙ��'Y?R�*b�H�F{���T�E���Jd�D60��<���҄g�۔.Y��@^m��D�>��k{c�Vus�����0L�
��d��<̊�7(w���thѝ�֑�cE�jx���W��5�79�I`>B_��}?�ʘ��	%�NB;�\dW%B�&��c* �z)䫳�B6�����m��Y��duo�C���
s3�~��'�y���0/���ZUJ�&�y��R�{��ˠZY�'̊.�X��>:8��	a��!H~D�8��f�l��Pǁҝ���ǃ2m�qI?ʮ�׫�Ї����C�_�=GE�Ti5�C���_� +�C�PT>9 ��(a������^#�U&zÍ3��.<��U�z���?�����'靋�h���Zm�AQ�RB]OC���.
�4�#����#�T��zԹ��V�k��4I��8s�7�>����J�Q�V��~r�=bެ���8!h$FxNtM����T+�HSV���D_���(����Ĵq(������"J��Q��_���\�-Z:@w���L&w<��\Q��q$���e��B�kv��N�=�_�����H���p[Y���p�t7�hϰ(��G����s`� (�e��+��?H��[
z .6o<dm����]���V�%��$��e��p�A@�����኏�`�Go*i�u-`�YI<������T�Ћ��Ma9WD�/9�3�r���jܒ�I\PA[��3#b�T�|J�K��W��,�&"�*3yr��Ǚt�8p�(�pk�Rq1��}������;��٘-�gB|k���̘��=Qޝb���hq�]1�X���w��c�[��W׃C�/G��~n[�.�h%ݑt�N�4@av����c�b��ky��!\���GO_[Pra��M���@:�e}]��6�f��J���V�p�n����cC4��3�Y���J�ۚ3 h���]� d�PB2!u@�h�AM�o�%�~�a�������.�^���n<1r�����������h�G��!,U6�����w}����� y��>��vI�@�I��$o'�����_���W���ڤ�55G�����G�LR�6��a������/u��E`c!��r�c�����p��t�S����5I��}��  %F"���`F;!a�>3#j�3n��+C��C���~C�
_oD�D1�'����PǛ��J��p�|�A�.�Y�� ��&Yx�$8M2��3�E� �,E���jgh�Wk�v��cBjR��H�L4L�"���f�KP\��$w��̸(M:�	�Izl{���E}��L��C��V!�������w=�}�L#�A���k^�1nk9�.(&�5��2 پ�z^r�d�`"�k���$�N̠��'��!K������w3a��~�T����U�%TExڈ��q)��Ӷ��ņz�Xv�WI�lZN�O=�ك_��n���N�Va1Aݔ��q0�mz�G �7XaB�������YIjP��&�6+�7�n��lFc�hr�?li�lm�r�ř�C&�D���t�\�w�XŬ��is�[���TTz��Hk�g%S��ʡ�b��n�o�0e�+&O�Jq�r#�vS��M�@�dH��핫��*���7��S������l둸?En��K#��M8&��I��s�b.}���+�o�\�V��]1�P{��Y���_dz�|�P����#����kb)F��Z�&�<g3�M;ٚI؁پ��c�h�g��(��j/���_����=��Bch��1em��H���Ze�&g];����2�8���YӉxhh7͵���9��7/�R��LϻKWۯ����>��a��(�����y�7ڭY
��ńӄ8������1��l
��Y���ov�fkTp� �B�_L<FPQ�Ga'�I���rf�����h,�d=���9��;G¶^���F���f���ɷ�Īx���6��VA�	sp�Y���s�0�c):�d�P!��0���\p5Q�`�͵^�%4X�Tb����̔���
'չ�O"��IfXڜ`�۠�ʔ�������_��\p�̀�\�g�� �����-���%���,��ǂ��?�v���+Q֯�����ϯ�����E�ZJ;�y��u��;;E�b���ҳ����`� �يk��\\����at�x)/�A��c!�e��� ��*{R�e�Z�^U�N����_��jL���lO����}w[���x@z����'-�WNZ�k���!V��Gbv�o���1�_����pl;|�G��-5=��WE���O���5�e胶�Y:a�gԍl������Q�hT#�N ��}��:�� z��DZ8���3�"I��V8�Z~�*��L��D~����>�`pL�t���EE��T�#_"� ���wS�#�m�(��X���+�V=t]/xM���*�t��>����We=	Ю.<���o�|���}a\<uB4J1#Y�E5�9E�rk��-ȗh�P�w�w�>=|�h
@�$`�Gu#�Q�A�PZaӏV����e��7>EK�<$ؘx��Fi�И��񺛏�<�n����f7Z��V�Ċ#��Vp/B�=�o� ���cɰ��^������?t��D��AN�C�[���AY�J�sX�/��Qb�5	G�\���#��{�(n����BČFZ240ҧ�;|z��4fӸGJ�Ӽ�BٱL�ݷ
v�r���k#EF��.?g�+��a�(��y�{iKa�Y~�ʣ��#�G���(Xs�JK��ҫl#�G���G����J:�兰���>/F���ڱ;��FF�{�r��x����k+�]z(=��*w�h@6>�e�������:�~�q/������
���{��p������B�Rύ0�N��ݚT:�AI}7`��RhI�)���׌�뺝�IΑ���Ĵ'�O�� �l��rL��'�z�a8^��G�ql��*�^U%p@:��mfE��xM؍�5~p�W�l@���Je�9V*&��}��"֎m�Iھ�*�r\Kd�^6�]b|����f���R �ݙl?��u�440���m����5�9��G2�X�i�u_��
�q������C�p��bq~/��6�s��	"��uO@�*��ǒ�"��dJ��{v?�j!9�����rm�JK/bْ�׹t�._��T~Q�#��R�A^��%�C��<��lr���V��D]�`=�U%��� 3K��_Qo�0���?��tt�����	���3�-R��jU���N��� ��"����h ��j��vb.�f�ۦ�Tq�b�l���h1V�)̎��+���hk��W}�d0�n�E|V��eu�X��M�H��/{��A/�
��@��!]��9�����gP�U=9�k����8�Z�J#������w������w����9h����"��=��C_}����쳸�S����b��"�{KH�lT;I��/���c����-���٭�wq_�� <=���)����sr�����.X�p}�Sha$ZY>V��-����I�X�bw�@�ө�&ݲ9�SY@���bƊj��ܗ��Y�X����'z]��t�h�i�8��������q�<t[ƽ�u�/S̺R0�!5#���Ll�;~ǎ�4ִ��'w����\Ry�E���i�0~�ncg�"�ߦ5*-��L|4J8g���TZ��+@�?#c@S���!���g���K"�<����E,��e������WMk�� ��ɋz4�K���
�f����Ќ�>=����S�n}6���$Y�?����&�5��d̢C�,cW%_S�}OX�Xف��?E�VH.fS
��3BРr�W�<`=凍�^�zx�f�6m�=�m�1]_r>F��G�K-<ܑ
��_�<$D���Zw���5s��o�9���r�D,*8��}�~ͱ��Ik=%�:�C�����$+�����u$S�ɳK ���ss��0���*K���}�6�?����G��LtǨ��1za�D-��;qC�D�2̻#\��8���I���g�`:Y k�l���o��l�V���$��M�+t7���ad��nΎ
�
U2b��SPY�����K�3{����݀��vR��>
�1P��&��S�$z��s��"�4��tE�җ$3�'�m�`\v� �}��Ī��l�:6"8�>]�<{��ϭ��.s]���~�%��f�*�I���`=Y�v�o�Cyl�C6b�J�G�kz�5j�w�� ��b6 W��m-���7�(������N Uu6P5�,� ���E���1Tͻ�[������u��j��!�6�e�Ns>:��[��@Ĝ{0Y-�C6��a�~��a��d�Ie�}�-�qF�b�֮%��������)�v�[�DܙXt��-�t��E���*����0�୧�ɯ.Sg #��&��k�5j#���jIk��9�
0З��j�H|��MFUEv�;�H-����v�ҁ�>�ho��KB5<��0o�o�I
��ӽ��W����v��o�<�I
\"E쇰��:�	O�*B�%[7���Bq7���
���ee�.�V�����"m7��l86�>�s��.��43�(pXn �}Q8tU�KQHJ����b�F峩���gT���5"�0꿲ʧ��8~��h�!.��"RXp��Ԁ	n`�zy��V�L[���J�u~';�@-��F�~�L�ɤpҦ��K�Z��QG��ґ�6N�ʐ�[�7@jI>
ͿQ��	�ù���LL��nW�DX�jsޫ�ce�e��W���Je�
�d\��8Q��������^���MQ/@� ����1���}ϋK������� ���ɶ��	e�5.�1�6[�B�}����mb0r�k�3�d�i<{%������$��]+��5�a�<��?w!�������9$������7윂8�k����';l �-�a�����P�>�NXCg����ݽo��I��2�B����C}n&�!z��V��O�cp�K��m�=��DHsݣ�cW�ԀCs�S��d�1I�̷�n�Җ�����z�)@أ�+`�f;�r��¼re�$0�g㱫 ����M�:7
])�Y��0ᱤ��3�H,�b�+��W�\�"0s1� �Q̪��uTi���`BR��K�8>�*�����뼻	i6�f����F����ջ���F�.�ٛ��N��dL
k�p��8�}2i���@�ȫ<H,���������D��]jI���1�(N���p��e��빙[7����N8L��s���p����ܱ� > �.���eH���>[̚H�p'�S$��/�c������uю���9ZZUQ��f98RzA���$�^��C@2��V�e�	����lnE6q��J����.���$�����n�J�t8{{�݀���?��GY;n"g]�&ӿ�]�p��vӕ�r�q�;e��L���+ڐ3�/���Vk��L����Hn:0�[��Z��Q=��%�����i�c����lϩ���>Ї�T��y�Q顊�d�,wظ��T���i�ǳ�b���q�=9\��7�N�|G�9۩9���dƓ�p�N�f���`����^�J:�<��Of�R�w*ğ=?�q�E��*�uf��d�+;�Q���ޫ%�:T���X<O"�f��-r��3Ҳ���%"CظWjX�o���|��9�w����!֩��� i0�j�?u��[_a9UD��&M��D�AC[gh5�: �����^[e��q��[�YJ�pz������]��w0M�Lv%�;I۔��1d�l)tV*��J�l{D	y�֋M�.�}��n5?k�X%LDY0��W;��c��!��2oL9�
�MF�qY���͇��㑍�:��x������/m��=������3VP $l����*Z�Fv�]����g��c�΃�t�D�d�j��!�r
yW��'��ޭ�d�/��B�v?�80��)3l%��G����[�.����A�&σΝ&�Vk�z�\n�nB�+N� ������s���3�#U���)���C��@�^YtV
>9oˌ.uX�hV��f�n���|�k;j�Ǘ�YS}]������]�P��~�X�Z"��$�ah��&w����
a��k�/ۙ�_
���=�a��@�U�Q��.	����C^.�C:}�G�IL`;��bፁ���q��ajn��)OX��Y�Ha4�v̼��ڴ��=�i4�>>N�[����B��i�g����=+b:S����O��h��n��U�mQ��cB'q�MųÀ�@��k~��D��{��'م������JnI�!��|Řܵ�g��6�^���F��A����{��j좶-�U��~�C܀y��l��=�NPfU#�[b����Ȃx�OQuQ��M��Pc2W֚��L/��j���>��E�k6\!O�//q��wA����@D��K8����9E�9��i��=���Y���49�Iq�O��+ۨd�C�#;� ޕ�J)`�d@��	Έ�<�ĀiJک'(� B�.�9%o(�Ø��d��2jH�j�"{>��cSN+�z�lG�;[.� �$%���aJ�_�L���X �V�NL$���_㨔�����K�l���e/WX�p���]��4ғ@6��-����p��3꾇 ��$�[z�~�P�pUK��Kj�TJ����!~�)��A�2`A�����sF�Ɖ��s�/X���K�Oި�~����qJ�R���c&s0@��UD>��6��]��LB�/T
kY>��M �hQ�NC�Ţ >i���\�Z�J>����%O,].�1���J��Y����5�����n�v�QS�Zv!n����O�,O�%Њ b�ɜ��;W��uhV�nc<H{c�n	!@��->)���1	�����H���v񬨃����
{r���2	����~B��dxq�{�,^,�������]+���v5��_'�3��[I*9=���:b�o�[�@dDФR�����>LY\#c��5��J r�bF���io�ǣQP΄�j�m��j]�7�����H���r�Y��e�5��p��6�3��!
����Cȝ������.a�)"e�h��h�X.SD��V��$A%!{a��y�M��d�J���Ҟ�qEpMY�W��oxŒa�>�� Ca�ֽ�l�8-�wa8��o*՝ԑE̓yuM��'��`�T�G�ZJFE����#,�آ[>�=&S��-J������s�M3 	w6 � N�x3yl���_� AZ$�5�uVHKJ�" ws? E���E��DFI	��g�C�y��@�mmf��N��<v[鎭����UYeY>��>�9M��	ң����%�Ģ��9��+�����wH*$:�3|�߼��e��_����>y�/~���κzO��P�>�OgQ����^	!� >A��d$�9I�͉�N۱WE���._��6eo���jQ.Bc+�Z�EG]Q�Dڐ*�2@��Dy_�a�+�
���簅[�DeS�s��a~�F��⸱�]�Y�~�rR��H�t(�,]�
���D��@�`�w���ږ#T�&��8����8���������$�n���*�<ΞKߗ��bwY��x��A�T����n�f��]�����_=��K(O!���
_�9��Ǧ
�L�g�!�������wpQ`������R��;��6�B5�� #٩4�R��,_ R� ]�,����R���A(]���b��ˁ��嶨�=�&N�bX�<~=�֙ߢˣ���Bs^Jn���AO!n�"�]���~�>�;�#�m7��������b+(N�W�'5�p�n��e�%�B�*��q*>�u{Z�Y���|����%��m�g���*�sβT\W�bke���S�V�ȼ	׎���l��w���nMP�}���/n���/�؁��y�|�y/�Iq�)y���%a'`P����r�(j(v,����0LRc�'a��> u���ݖ�A%6��D<$�7�M��#>(���b��e������Q
�� �����̰Mu���xDV膩�lf��>[cG��V���_&���R.{]���(=n�Y��ۮ(�m`�6���ߪ���a�0/c� �=w[������)�%�J��`�� ;ы�KK@?�1-�9�ٺt�ķڠw������$�~,�������JN���>�V]���Uʩ$�6�FQ�-�Hf�������~m��i^ �̴?h`� 3���/��#R��{\Q��φ���j6㆒E}d�	�7�{�yL56ntʒO�J���穹c8yqrx\�ZI-뮆O8���$c���t,�O���wdS�
]�M�*�!:� ��Iaa�&]�Z����kR�� �e�����e��J��	h�9 �y���Ɛ��A�}��$�?>V'gm�������X�*t�j��y�O��^Z�Æ�x������M�G���_M��eOC���7ܼa"<ԡ����\�H�-:��^�C�4����п�C���x��Vf��5���z�����7�<���k�����,_�K?}(��"X��әZ~�ehw'{:�ݍ"y2��VN���亪����1G���pf��0�=���0F�nQ���a�27�GR�?�`8�BV�60�C�;�cm15j�Trk4��i�z%:�&D̽��R���s��P%�Qq��{�kꦖ���Ճ���֭w������DJ7�γm.e�2@����l���r�h:�*��z��!?��7��f`����Y��3�Ͼ��R�h@��S��W>���Y��>���i<���e��k;�a0BB�ቡpn)q���㛁�ÍT���s�=v/��/�3[�{��'	<w��9b�� L�!�XI��&�?ӵ;��ѠWޖ���l��,Ӎ]���m��)77ÿA�8v u9�;����Y�ɛ;Oͮy�2jD���v���r'I��Lh��Q|^�HH�b�Jp�	k\ZB�ϻ��3����;h���;�>�����X�T],Iܱ��U��]���f��p��^s�Q���x�F�=:��M>�������=��,�*k��7*�����i�CB���skZ%�m�l5����, �-�ҁe`�Mlؐ��\�F5<�ٜpwy�n���LC�$S2�x��+�a:�����F�!�e�MH:h�}l������Z��!}Ӷ.LN�(�$��]:6�<S9VOm�����Ѭ��$�V�P=F��]��Q�s�k��;�y#^(oj��;����-7ma�/��$_B�.�ky���E�gu�p�p��:xi�Ep�й���ayl(8�"�{uA�R���Q�Y:�)ų��F�Pݣ�(�K��^� �/Qь2#�<���i�^�^i�V���p�Ug���V�V8�F�i��<|o֦j��ε+w:��/Ŋ��t4�7���)�%�g�4ipWg2��͢P�i�>�܈�XGn9���C.�.���R��y�~d�癠6�F�q0�DR;��_3�	b(�7?�����=!�& '��6�N�lۀa���7�
���0PWqfo�BG�������!=r�,5~��qLT�吵�v.&m�vI&E���M=-r%������<Bm��3Fѵ��J1\Dg�N�.�Bk�Y+}�x.��|0�.��kK�;�u����_Z�� ��F�L>0���yO;k�p�������h�z�8�ژ�� >���z�]�L�+��`�??bb�lT��S�
�\�?�J���d�+jqԘ����t�0� v��t�"u�H����ی82�Bi��Q�T�GBep�FZ������g�qc�3�.���:��Lz	��OУy���_��ma��?K4�c�QC���z�b?V� �s�zD7���Ŏ`��8[���LF�6�eʢ��D��D�y������*W��ʟP��-��%�<y.�J#8���0�R~�Э�������c(����s������T�2 =s}!�Y,p�_���u�n�
��MG�k�{*<���y}�XP��Y�8|��L	�"q� cF��M��N�XA���W�2�է@�!iW�4�=l�����}�#�7�Zq��e{U�R2����GܔH?�h��ߕa�5�� �jN��it'is	洷�m����@��xf�Q�,G����[O��\�fHB�8[�x�;�g���&\<L�|J��i�c���fc���8� ����l�2F.i��jqW�KI8�h=��	g�����
sM�"p}��M��F�0`�҉1��w"5hm#U��~G���cކ�v������>5IX�g^U=��4{��Ϧ�z�׍�)�	�7.q����C-��+Ȯ�H�����M�SI�U8�^S�e�{�({d(`�I$F*����9@|�䨂�.������ihK2�A���VHc�P� ��+z��;�K��_3e�w�v�]2�-U�6�g�Ћ����@������,��x����,pd�	D���X���C��9X\D�b�?)���S!Ԍ3�c����2b��#/�y�k�~X������ݚ+QRu���;�jZ�x[W#��L��1xV����I�E���·�")cs\&��R�� ��k��cU�Ox�掿G�)�O�0�ΩX�x�bRʍNCm��fmt�ƺ����a�1�Z��$�G���p=�o4F��Ջ���
z�� �R9�tŗ�/�'�h]�I�W��5���m{��/����M���>�o����,�z��>�#eIaY/OשSXr+C!X�%������1�lG�{K�콁�E��K�h�-�no�UW5p=�Iv�X�ը���*%~��֬j�h,�����h�����'J/!�\�ذ&~�s:y� ��E��� �u��ȋ�ӧ;k��&h���E�(�+R�U�j!|㺝g������dڵ*�;9L���gZ;E4��ſ�t���,�&x;BF�@]� g3 Fō0�d;i�J%�~"O%��{��8X��!��ejd1X� 긅�|�� es�;��'P�H�Y���2M�ױ�	���t�b�0Ek�+�#0�ʠwb;�A�@<͂�26���<�'\k���z���!�ơ,m�����Y�@������b\�'SY���>�brg�7��,�2��{@�{gLʹ}�7'g{_�I�E�l�y��&�[�գ�l���3�d�X����Q
���itW��8$�-ZPǹ� [�<A�E�����Ө;\��'�Q6|��lv��F|�w�G`u�a2��!3������N���lL���jeo/���kkĉC{��+ρ�Mk��B�+F��&r�c�ƙu����a�CY���z�Y�v��W)F���v�2S�N4!cp��I�M����+�N��vy9>��)��H���: A��0��;����X�l���I�6%cz;f:�5�_S��ɞQ꫑���r�K��_�)eھ��wy����6p4�'�R(,��
��v~o�"�m1М�!���������w�����7'����M����h�T��O�M&'�/I��@���=@j��J�a���|z��,�g���$����9��𩾱��ޜ.��͙�R|:�q �1X�oTܴ��~�`��q�����9�8/��\�9Jsz!�ZF^4��]_�H���W,�W>�{�Cs6��6lp�R��(S�� �Rx��[�����4
��jH��7O��`}�Gy)Ϣ�4�	r�R�����ѻqk׉���L�5�j���g�[JK/��_oC�u��3��l��e����;�LQ:�%QD���������V��򼶻p�)ē������) �Sxass�8�p6C�{��d�#m���|�E�H+�vT\��v�Մ��q^ay�B�j��ξ�e�=�+;�|_é$��0�x�fgR"w��-���7�P'�_*+ϛC�.ȑr�o kB�G�Ğ���_�Ö ���\ܘ�M����F\J)6/n���>�U��{�λ�8���D���K.����z�ɒ�Ė�Ł�����V�_���?�#�Ե�{^����V
1n�:61c�h3�O�=�t��Y���3�k�U�Y,nB�P�=������K4
w�*�Ak�T���8mk��	��M�:�3KԻQ���I$�~���&
�	�A�qJ����d�rsmg���7�LZ��k�n�+��Iŋ\����ʵa?�}�
��i�ͮń����c�W���GK5������25�G��,�)��_N���="V˻��f]Qt�B!�Cngk��"^:'w�	Z����;��JE��J[ߐ��%���;��&F,��x_E4���/Z���~Ա,�)8U�.��i�]�3����/BU�ck2<��m��Z�LKʸ~V���+[]��=�k@x�P���`{�\�*����$}���Ak�7�Ƙ �a1ߠ�Ǡ���hMS��U6�ub�q���;�^ƺ�G�{�@�\,�h��`M�P������$C�!t��Q!���W�/�/�6�]��j��5��1��	Y�����Յ[��	��,m9<�*8d�bÏu-ĩ\v�X�U�Љ5���Dh�	(*�#N^�:���ʃ�[;�#;���z3��Jޮ�%M,���/e(Q���Y�^�~-*:Q�����î�d|l�\f{TY:\�?{��w�Ц�z L��F�	c�g��G�7<��,�uH�Ba􏩰ң��9�'�}=x�*I;K�i���[�ԫ9��|��>�{��E��^b�}"28�/�;�9�n4DR���	��h�0F$�g��O1��.9"f�8��H��!����L���_�[{OΑh��<���T�&٫P�V4�bME��r����v���ʪ{-V��?��ME��:����b��o�w��5���<�a�ٍ��zĕ/��7�xF#��B��:��@��jE�=x�!�y����:�
7�(nmM���">�_v���q�8e�����6ȡ�����%&Q��A4�܀�]�<'e�*���p+�1I�S�f`A�"ղ1b�9k۠>����a��xa.�s�!x�c�MĈ��������@|=|����t�)m��iW��+�����7]la�\g<}#����}�]�hc���eƎ0.�|f���*�)�{�8\��j}8��rz\	X��.�dI����3���������?ML{٠�N޽_ނ�9�=5Q�	����e�b̻xQ�F.�D��`������Dum�O{
���!�by��Ű�3%>��Xo�g�0Er ��#%9�P�$
wU�d�#�l'Q�Sw�s�I`o=6�]HQ�WQI����"rP1�Z�>�׻#i��0��Z�V�<\=3UoB���9G"�5UF'G��p���s�[; ����;�Ȑ�(݆�<躑� ���I?L�$������l4a�
x��9@W�?�:��}S���7��~��2���=����y#�;3���`��iwt���跣}��[�))$�d���t�-�Œ����q�V
7/�鿛u�*��:��n�J~z);�� `�:>��mZ�UIY�UF�cK��؎���?���׶����=|ަלj�V�1����f�`�z v�8�8-e]ĭ��2��k������G��~�;S��3���QT����*%��Κ�N4�NS?����]!��ɬl�pp�(:/4��ǽ؏�e#t���%^���N����*��@��m����Ql�Um��~&Y.�)����_�"`~��/�D~2�X~̩����q�R}�X,9|K�q�����;�[�T��qʨA����A���Q�U&2?S4�Q���Я����f[�5�#Q_7z��)i�Af�x� ]JC9�m��	��Z��r��[��@�ϑ�J�HNk1�UO �%3�o�l3�B���-���Y�#�8e�qtCc��`J�c��~⒀���0�����mA�5�I1��)Iɘr�#)3�*�+FK\���,��r-6�^�8Ʋ6�n2ߏu<w�吏^�^0�1s$���y��oJ �F��xU�H�O_�q�J���$���Fk��r�:��}���	!ر�)�	�i����}�֡�T�68m���G�� =h��}�E���vI3Yp��Ĥc�˙ǗO(�y�m�h5�z�w�p����^L�{
S�6�aaݶEy���|eq1��L��&+��-�.DM��gL�!,����W5T�ty���J��%IQdV��B�҆]b��:�ux��{���>���F�0Y��i,�I@�q��/:5I������V�����M�ޙԉ0Z�#�W�h^/�E�k�Q���0��.(���!PdS�w_/����R�<Y�<.�7LEc~�E"4�xV�W ���pţ�{���S�a�W��RO��&�F�����ş������5�?��]�뺣Jo��|���n�hŽ�����#�A�Ҧ���n��wտ���Z��w��nuCJ�ݗ`P�SS��l��Q�sT�GS2�����B��16cBA�;�f��ܾ�ԁ�I�7S�[!
C(4��2pʘ�2(�i���t
uS���d\�j{GZ�q)4��^u�X��(i����*TWQ�y�w]�7Ñ��lRG��;}NU&U�G8k8���Rt��ez56�.;&D\�c"��9��mgR+\>��|�/��n��t���_�պ�s�����V�t��@$I�!��Ab���_~?��B
�v�i9�9Y�?�H�^�¯�A���>�9���x!�S�d��zj�c�����̻Y�c�q���!�x��m�Pi�߀�KC)���H�|6b�'��q�#�oO �t�R?�xe꒹�@k�ұ���3	Ȋ�/���!�in+.
VT���x�Nm��¤�J��D���8��'�i�������fl��Og�QRC�C�*����'\��O�6w?��.�&��ʇr��[5Q�1�tE�q���߃9�ݮ���pv�ה�H����T+�Ѕ,�NU����̱-��#���]��r���Z��p����L�ܟE<ڳp7�w�	���P��Q��3!�hC����@��V�G!Fh�����lT��&�l�<U�Ѷ�ff%�k۹j��� ;ʯdB$�ym��'I_���y �q�VY��9!~�{���I��X�����&w�Z��mH9vV{��?�� :����5fk�1�&���7S&v|´z�Pl#��-��_��&��e6v�w�A7�p��{|��0Sgss@�4�0&�̾�ݩ����Y���A�-N}�V'^��g ��1Ub:�+�CdUO; =~�ʱ������H,��� ��}u�- ����Qq,K����� } h���*'�p��x�P��Tu�s�xM���g/�����20��߼%�X�}~65;c����#0$V�%�y@[�<�Z�G:OX����J,0���HY�,��>�]��]蜛#��<��I!`<>���>�v��
����rk����8���=|�*P�R�^5�A[���Њ��bQb�Q��F�DTUZ�&�$��F�ĝ,u�eخj�����o��'����n�T��
��- �X~�^�&�OU�����VI�_��VUY����~P
P�.�e��!�R�3���X��^ҀV�?�M�h~?��}�ǰ,�����ʚ�_y0@�i�x:��+�>��v~��,cq���c�;�i�62kJ�L����S�x�xv�ko�Ty�;��S�¤��p:��U �Ln�c�;$.�3i v�dV�	5�YD#<�R��[ �/�*�[dY���S6��$�3���j0E�S�®�A�k�n`�T�n'6*//T�c�s���&�F�����]�>�dcG�e�Pʥ>.����7�Y���������&ty�V_�j��6�v:
�an�{=n�E���i�c��U�d�ʃc~��x��ݱ�O��aN��(�{�v�D���z��f�Tڈ&���7-�"]L�5�� ��u�k��k�.�*�v�/RL��bV���(A�7��pv�"*B������ K��b�6gn�&�����cG.p�c��G���yh�ה�	��1��s��ih� ��X�$ٌ"z��z�Or.�%�@g�PRFV,�'ڗ�Ak�=�L�A宸���y��,�ST��X1%���6�Yv'�Ow�9 ���{#��:v��+�ϸj$�,�bhZؐ�p����#��ј�m0���d�29���ѵ�R�Π�[S�1�Y��}<6��<��x���_%�o�b�ɧ���m��A
YC�P����[����t}��w`� ,s�#�������A?���I�\��]R�w6X���	��ʝo���7)9�ϼ��m�#�I����7V_�>����O�������::�F/��
2����+���ud���:�W �u�`doP朄����kd"ܢ�h�(?:/�uzc���˰�H � U`#zS�J��Y^�f������;�/�������;��j�5���?A"
�ʄc|D�+	��0�r�:3l��A���/�o
��)ya�+Vr����Ki;Z֙|�QS��|:�n�^��Q��SXV�W�A�W��/Q-���=��,ϭ��;�S������\G{��r`b_���/A嬂KpR���<���
4��spИbI�4q�)��S�b��'�tm�i�V����Oct�i��<����������d�<�N���)���(�?f�X3��4sG��I~Q%��It��	�)v$�9aa�83WP�l��2�)��Y\�J�dHcH�.�����Q.(��6GУ<>>�L c��}c���# �'��
�35�T�ԁc��f',�32r�������fxH�9r�p����z�&�599p���@�q��:�m�o'b����ޑ�_l�tK��[r�Fq9:5"��U������2n;���ѧUThӃD��3�6ka��L�;�zO�$0ԃv-�0���y	�re�z��cH�?Dm������O��#�UtӐ\vӉ���c��I��XcX!�:a�L���߸��ʇ�@��>z�@�zqo�ay��l�M�13S�"��6�*q��*� �i}���)B�����x_�b�A*2e�w̃����m4����Y�~�s4��^�L簬�UILQ�`U}�x��-��Gp(8���虘x!����� ���:$��=��"�3� �Q2�l��	R����7�2UH�cտ���U��#����]�9�mV�Ĝ�/�T��k���(`�D���*�g�Q��af{=p�N_�S�.�"����*n���"S��H�Ǩeo����I�A����_�\��F6D�r�5����Q��K�>Y�W!����|�|���@sI֧�o|Q\c��-]"Px1�:�Yw;�����Ԙ�#�i�k��4��g}"�@�Mp	!�p��c�4��qS
z6�]g�#��- �w�d�n�O-��a�����o���;d"�InQ&%�>%�b�ϓ��A��83����2��2��U�|��[r�߉�m�N� #��J�m�3�3���I�.�C`�Ѝ�2x�f��4�TДbs�5��k�oL�UC�ӕ_��v����A>��Vv�W\��l�����n&&˨3��I6ۋ;K�M�=�	fdK�!�l��*+�<9�O[��4 $_�7���b��Q��sqߢ>B��tj˰8647=b��]U�V
߃'����"[��y� �M����!:������#�Ф��Q�ۏ���4�M i��_b�,�C��ں�ˮE.<���	_��+�S�.6�F�\5;(u���&��;�%2�\����<ɱ�1�)�vX�����?��KG�y��(+�䑓��	@x �}F ���:|�C��aԤU�lx��J{��?��;�_O�����Z3�--�T�� ^DzD�	�I�+�j4^�}~x��@�]>�e\���Ul�;2B)�/5ǥ�}l8s�8�%�v�߂��R��N2ʔ��E�^���F1��8�G�ß5on��<��h��^�&E��=�plG��[�f�Z5�4�A/E���P����y�����>��[��J�f��"~�'O�d��TV���cu{~��KՁN<����i=x��m��/���:*�+�ەIT��ˑ��oO�]�^�r�ȯ�A��b���ٲ�a9���l?e��:�ޅ���O����maj;�okD������Ƒ�_N����4�����ʕ��VoPs��-m�i��dZ�6���ζ�G��`J�1�^7�1�vPM��璗G��E�6Z��&Y��2���R�X�1����Cc�D�DUu�>R۾�E�����"h~.A�	U�
�\�!���qIY�	-~G�P���s��Q�����۵)�F�����H?Xa,Z�^�ʳ1��2�*�!���#Ř{�v Ȃ�@P��{��TӺ�
��u^��b�Ή����2�>�Wt��K@�H�`�]�^7��:�_gx,+ZK�e�8�)�%���c��
��@P��L}����Ns�#��{�H�t
�7~�AU#� �`r�P�9�&��s�+67Bd1}c��� t;��,��bh�EP���6�-!�AE�qvz�zϚ�$_��x�AxJ�v��~[�\#Ö>�a�R$?$bgt,��i3:���`�I�N7�8w�t��b�_����}�;H*i6!� m1��S���-����A�C�m\	U�g��9'"g�-��Ɲ0���n���6;߲%K0��[L��va�	sv8�8-��-z�4mw�J�{K�SKg�Xn�=$?��w%�t!G5C�P|8�I���q�K������ѷ��}��-�h5����kP{��E�'��iVS��jg�$5�F!��n��鿃�	��ɘ���Jo��	��J�]<���3��6*�$癯�567:�O�26�6Y�{]��k�Vj;�m\�[�R��v�a��Q�'�U���*5��dmb�'��i��F� =� �oY`�z�TQ_.� �x��qi
�B!�[��:?�5�h���b��7A�M���f�O�zC���*�����n�W��긍Gjɰ}ZX1$�J����$q��Y����+5AZ�IL��1d�yx7"�.M���`㔓�{:�sQrC�>訍����=�FdOn��"��w6��v3q����e:�(k:\�2���k��M��J
e�`x6�|�$�G0�`׭����w,ljt�����$<��q&~�m�/���\��:> ��hH��i��[ｅ�W\�#�֯U0h^���]v��o�����&ŵX��dŲ�}���"(T�	�{�Bd�疏��D�9 ���C��Ky�ͪ��,��=RGˊ�W��%�F��T3X��~�̲��ę���0�l	���gF=�J��N����a/<�L\�pݪ��A�.����;�p�)�xup~8r��=�2ͻ���j��q�?4�o/J/b��Yo�+��E5~�O�d�nm��*[#b�+;e,	�¹���BS�E�\9�F-����ԡ��:5$q��&Or�-*�R?�E��3����J[�3����G�.�-�/P�a��k����j���qEHԕ�F�Cf���R�ަW����C�f�A�5�L��SU��3]a'_�g~������i�w&%��Hp��W6g=���Ƶ�	���b�5��%'�&nـD`Z�y�`�e���?��J6͸6�u��*�jL���&V�F��m2�"%��+>! ^&e��m@M����Az���_��#}��#%76<Ei�����R3���խ
�Q�y�[�~C�A.��$hCь��&KtUi���c������Ŀ6��a��bHȷ�	 ��>V�ld��~���-��0�D'���i�����_�z��j�,�<�������{�	��|�ೕF��e&�<�J׌�/n; �^���nk՘��e��e�ۍf����B�0�ϡ ~2�u��+A�B�4�r����7p����q��;�L�|=MXPblff�����$D�[N�N(�'�\R��H�������zu<�p2i�S%$
�"`'�u ,,W���Ss��L����u� 0�.g�9ͨ��w�*�����̛���odA]��<eb[�F��*&NB.*iܾ�����)�Ò��uĸ	$J͢wі~�&, 4��N���6���{\;���� �����"�x�[>�k���!s�K��&5E�-�%���g�Y�W/ 1���#\�yc�\,�x�s)zgdM.��?BKQ�(��\..<�S�I�C�W�h0�ڷ�� �����!"�c�x�y9y�::��qD`m�m�!�Y�L���)�7O)v��?�ym�{e�y�u�gb���tJ�KD"3~�,.69e(��@ܬP������r��ג�M�$H�m��R��mF-�^��u�W��k��Rv�(�	��Az�Uv@�D�ک��Wc-��E�t�/�i����,LK��BJc==�.��UN3�ߓ
�٨�>�a��p���M��'U�M�iR�5����4=�~�)c���=q_>HVe��Ƴ�,�tH�6]@a?Yl�)axRr��tP2 iH�+Q��"s� ��$���+��?<��>,��Υ��'���5���y�A��w��.��`a0�/���2���ç�����S`�)��N�dW���:���~C!p�*��P��F�I۫�)Mʸ�����p��c�x}��������˟"��1�}v6u������=��!F�-��{b2'#���Ĉ��!x�>��%�g�?WrD����1k��$Q��:=��h�-yYJ#�z����P܊ v<-ǧ��6p�R n]ĵX������]�V&��Fe[��C�	�C6B
�w� �K�hh�x�EH`�ںŜ���˒EI�s��-|�,�B�Z�h�˛S$\ڨQ�|�����.�U�@��$7KU,k�6��L����Z��������f"�S�>��"�ť�����֓����p*�~��/#.�0^f8L��ê��!�ؗ�;�^��vRY���W{��?�9��̀[�����0=�`_���+'R�Y�9ZϜ�0�$��b�L�I�dw�E�L/ �I��B~��#�C���G������gϴ n�8��o��)��nM�稄��&[�IF����d�f� ��qd�u`�EV{R�f�it��5��$l1�-�
�`�sX<HVxG���}�lWmV+�.Ho�N�����^��
ۋ�Z� �o^�	1o`�t�1���m�7���f�jr�F"��T�$?��M���<��(���r�:}X�����9��*��Y~�3�H�0�	Ф����4�����?�Z6[(G ���t#�Ù"�����Cd7�D��gd�-��G>q�H=���� ���ֿ"}"�4nRa#�/+��:���**l�ާ�����1s4H��%Tm��-���֣��T0"yh ��n/.�cd>�d��oMI���nO�ۂ�aFh&��o�h!��ہS,�FJY"�qu��h:Z���?�e�~	^�h
2���xjW&�b�.A�$֜��$FH.0Cn�ְ��B��Vn����&����S`|�_6���H�R�	P/$�s�r<ӳ�Y�}���B?^.�T~v)9�Ć�2`���9�́q6n��ћ�fB� 3}'�����4�x	~zpu���� W��`p6"bcQ�<�s�X���0膴�-F1�B*�'ʙ��w�rju�]/�͜�6p@�юCv�!g����w��x�4�~�������5�R��2�E�ІZ%SrC9�)��朒�����/C����<f�V�H��k?�a���yK��p�y���z���x�R�J[c@�_����:�����2\�F�y����e�J]�h(�0����{z��W��_lq�/R�X>����hSۚ�C$���2eA(`rp�T�m����k��r��*p���4�j�������c�`M����^�(�g@��-���M���{���R)���3�?����1{ ��x(pV�1S[���"��,Ӭ,=��OߟV}��%W�$�5�p�3�b�����r�%��I٨��^(�M@��T&㖰�6���!���\cn_�X�L�R)a� �	kc��p��	ȳ}�j���'d"����{�+	�vF�b^h������W�T$��b�� }aW��$�Q@���� �Tߺ&D�߰��[��0+��Z
��uB�W/�C��p�Pp� �\d����P�ś>���X��~�jQ2a{�p�)�"J1g�7	.���p}�1�v;�LJ6�r�7��A���த&L�)���}�s����L��)x%��
�Z�����P
�槞�g��_�y���S:Yb�
���x�2Oz��q�A��5����C����Ƹ�\cj^P�}vp��. hp�̲�(������ܮe��L��p�ǭ�7l�kJ�F��EڍT�����_=�zu�\���(��h�ߙA/&�2�I1�~����Ht�cH����H�`�N&GY33�Wn�Z_Cuޮ�����)̤������u�ۖ���M�p>��a�	;!&+��
�	di�0f��	y�t�Ӏ�N���*�5�[F5��+�8�1��wo�~����c�bE�q�F/�:�~����-{4S.Ҩ����L�Ob��ȝ��2�n�'�����ۇ��{��я�
rR��HV-^e�Qu�������C�e�S��I��{ڔ9},:��>�%��-�U�F�f���6���~-Ǻ�q��2�D�8^
�~���2kI�:ұ��\�� �r��'�v��	_�>R�9,܆;���g	H��g����9
���S�W������D�&�Ts�c)�A�矝�H�!'�8�������gf[,�B���|g���1�\47�QƆcPޢ��X�d��p�ۢ�`ߒ�SM[8mTi{q��!��_����ݡ���Sk�/O���c�2)�� }��g�̷	�~�Ex�G�>@5�Ni�%�Cd]@�B�GA9����Q�3՘44Ni��Ѵj���:�w�,���
�T8�TH��w1�{��F>��b1�þ����|o:��"��@ҼÁ��P6j�k�K?�q޺h�P/���勹Lc۸h?�䧥[��b���������ϓj�>���ʯ}c
_k�"����U2��&J7������/M�ij�̰h��#U5i��z��.�E���ww�����Ō�����٠��o�9�6WY�PV��&���*�k���I/���
CgDvy�E=�$msZ��3���S@8��ޮ,?uS�nڮE�=z�Y0���p@ּá��SK,<{�zx�]Z�����>=�H�0Y>�܀�xK�}��1|(�.�F~.�D�)��@mEF�b�\�]Y�]��7$�z�Z(�̳�Qʳ�h��������b��<]+:�����c���`!h�K{����%Z���+<#	����;X���z�W�'�K���a�sd2?��V*��a�W�G��~�MEѸ�t�����#|���W���I��[�e�z� d��^�$&>�-�T��C���k����L�	����9���&�Jo߅<�F�ef�ƹ���n1�ȁL9?���L�
��q�a�2��\�{�e58�nL�{�����֠ha�;f�y7�5F1ʩ�DP�6�����w	O��s��G$H�}�G�с��T��8 ��s�5�{�\���s���*��ζT|����Y���!9?-Hh�����q�F���`?Dl�"�q�-���_���v�2� �L�U�v"�]���#�6���Q϶��0F��03���� ����3��8VC����*}.s�Q2�DK��ъ��k��^���E�yK@���g��(MG�(��uA]ܸN
 ṇ<m�I�7%W%Ìam7�'���fl%������BV4۲�t3�e������58Pɸ�iH�!$�X�{Zb={�f�L�׀(nCsS&g��K��l�E��b�L��B|�@�������7CB���,`��Y�t�U5�t�+j�Qѭ��pb� =8ӹ�&�ˤ���5 �@�3E��Q��H����� ���w捛O}�-"��RN��q��{G�~�
:U��8_{B����r����k݄yg��s�����|K��+�nL��V][K�Ѫĕ�I� �t�@O�WYoqRZ��$�zoMd1��`�������H۟9Bo�GiO?�#s���R��v�пKa��tpE���ˌm���X=��W��T��{� ��o\��:c�����NiOq(�̀������G�p
��,�=#`QS��B	��+����Y� �/Va��4�Ģ!���?,��`D��Du�~�C�A���|�D�K��G$��-7��_��3]�`S�nҙcΓ�5�CH�a�����Ktx_t1�)��e*��4�O"b�ѧC�p;G�m�������{`�m�8��]M�B1Kj,�m^�F�*t�^�/uM�Y�[��B��xaFXbt�5x��JLI{BH�J;����H~�j��~�7ש �`4~��^r
Y�W�OPD	X��{��3_g�C*%��v7�Āù������5�/�ג�m�7$����Q�pDI��R�{���a�^"�JE.�a�!�I���$)Au��t�A�gA�\,������dQAWaܺ����������$eq�y.Y��n���l�:�<�_�Վh�a� ��v�=3�K�v�W_��~�	#\�r�h��L�#�<G�A�V����i�g���ُ+�Snw;�s�!�UL4��{�Ma� ŷ�v�D'�=��)U�*P�ƞx
�^���M]yr�@���/�ICM2Ρ�Ɂi'���1�Y'{j!�y��C-T:�"�FYY���f���k�������Y3��5��3g�2�0��|�B�\�i�N�#�a����Pm�h9�Ҿto���@f&!1p�!��K��dV�i�R���!��J�K��(����M$���wN�׊����7��v`Ċuu���l�9ct �1��{�!��q!�&,uOI$GB���uW!��PWrm�5�:֗��������(ly����G�k�)��SVab}���NY8{U�)j|�����|��j*�����E�!y9OU�U1@qŗ��p.�D�G��+��I�V��9]��*5����Z�k��F�_
w� �A{�+�ʰ|5��t��2�$�o�<��JPeB���5�b�`�@��>����JeV	X��f��V� nr`���ˈ~��v�6�n(c�����)g�XE�I��3*�s���A}�0�D�@gr1Kò�S L�BS��%@��a����>J�����RE�\�F�s�p���g��D�Ĵa�vM�n�V^[�]����K���no��Q��i�!��862<ԙ)V�G�N@a�ܯ%��et��@<�wa�@~"J{�bJX���*v6Z�N���5]�Q>qn��|��\`1��X1���\�"���mֹ��ƨ��"C'Ӂ�3�0��#zξ!,)��> ,&�Z�tl�.� ��.W��t�|��3Ҙˮz�=旤����)�)U�"��vo���҃9٦�Z罀*m�Ť�+ɇ��j��Ã������'��T�6 ���H��K5��;񳃷��t��+�a�L!t�/8��Q�UT�C��nd�[�%��MR#JҟI��'�"�o[�9�5Ƭ3�Su輆L������M�YaUd�-osG�ٝ�rkߓj��� HF8A�]���m)�����P���E1�S�G�Y`�@x�"����i&."M�
�C%>� D�~�R��8`��*�QG9��a�F
���l_���-�핿��	B��a�<���&ʬܾ��`:���T���D¢�"����ؤ��$|փ�-�h_�?�������Re�)*�moV���e�c�j�(�]Rߒ�JY�'
o�h��ie�+!乕���[�c��R�L R�*d�N������X��.&2e���-��A��Je�y��9/KQ~	O'�CY��	��ۥ�a˿B.{�i�.
g���4����G��z�Ԑ�v5�̳�����E�?H[ �5*Q�kzń�[��M�{J�#���7(��NC���f
�4[������-d\QW��fQ�Pf6��y�"9��n��w��`u%�إ�(f�=��'���ȴȽ�h������� �F�L/��V�L���C��A
�Iq�V*E0��~���^����.�qZ�?��`�^z���058�OW����)�NpD����څ�}SHwj��O���m�����Z�n�:�MY����Ղv�cF�Z�ly`��僡��_�
��9U��yz#Quژs8{�{�<("�i�t��_k2�`��t5��Ɍ�V�F�!Ca�I�8�{�Q���'.�l�Q̌�ܫ����n�X>M˪'򱰲2��5Mw08�,��}F~{_���->�O�9�Qyᐖ�3�3��	�4�<��j�a[|�_�ͯfʒ�J��إo���B�	nA��y�;=�:G�K�d[tn;U��^�z��5��P�I`u��ʳ�����W�>�8�uӮ7X;s��<�ڑ	��!��=�Tyі�l��Y{UŜ�	��G:*��k�uX�-G�0��{`t�J�UOY��ԫ�z��=��f� �8l<�D�<���*6X���Z�Vz���@=�Y����ӛ`i��g�|힁z ���+~,�&���EՇC� �J��`}�	��áK$l��F��n�׷�N(�Z̈́�f+�^s��B�=�80yC|��NŇKB��4o�����7�Al�k��k�F�������O�F�
�:J����gÈ[�h�?��ݷ�ҡ���i�!w	�E��u�<��s�(�	aH�7��b���[2 �6�&��_? ��R�1��툯UF<�<G^%������GL bp,.g�Z\����]��>ېW=�U�W�7v]Y�W�)�o��&%�f�ʬ�<-��>O���MNN�J$Ni|:�6��-�D]��z��p��@��q��u���w(B�:M����;�\�k���;3a O�3N��l.��Sg�0���ȧ}H� "'0�2ytaX����u~���8����G�c\}��c/���uw��/�z���zW!W���_���n�ڹW�|��+�L������c�eV���a���r����f:[���3���:,�&s 2�չ�t_�^�	��Ņ=B��1Z����4�E���9�S3�5���'��� >�h��&\������9����?�}[绪��n��X�D�<�-PFi��7����l�BHe���Ȓ��	��r�`X<ls6PxA��M�u���rRѺ�@"�_�[m "�V{�]�)�#�Oɤ���Y�{U:
ev�_�臱��J�O�0���7�� �5�fTMy_R]�7��jm��n����Y��z�qE���r�� Z{���NL��ܓ1����"�e���(+4Y�=�/��6?J
Ay�!6��T!�]��Ma�	;���Mƌ���ԑ�g�p��
U�O!c)ET$�.b0����ԋS�%�[K��C��X�svn_e�C�E������e!���
)]�S�n��3��LV��_�*�]�����_�pUt���SgE'A����Z�?�
���ʈ+z�v�-��l�TW)`.������ռ�ۚ1�=�v�֠Swq�/�o(N3`rM�'ݔ��@aخ�j\��������n�ct��9p�j@#��E�#��)�uSO]�`�X�jz�hm�m������o8�i�X�!����P[QJ"3���/>0����L ���Տ��cd��`�q�|O���5�9��R+��o=�ҝp�""����ٻ�$�F�����韐1G(靹���QA��4o�j���UhZVy�c�A0MO������q���_��9��9�${�S&�%�8_�H=_.�%�����7��xߒ�/���6��p�hi�"ހ��?��L�؟��{{��#AO��
���|������kEHx)4� ����祐n�;杰Fg��f�=�Q�-6��Z�*�*f�J�,M��듙��((j���@�����pw:w��W�����&9����E�a��wS��Jd�8�z#S�k8�*�N��~F.���-'핵O���':�UFy�N��/�Ǆ��$��;��O���?���x.Y�~��e�эK�σW���LD�$1Ou���Dd��� D&6nw�KO�7A��Gr\�'^��rM�uҳ�R#gD�Ļ��<��b��mXrQ���S��N?��Z�JF�h���q���tuQ�C>���oR� ��Dҳ֟��D]�+ڹi��vE�.B�Glk�NWl�Ls����{"L�׸M
��Z�]b��������2I垖���4]헗����@�S�4é��Oq"nj	�n��`n`>�=�z:Jg7�L=��*Kl�m��:�gk��ƙA0C[�>���Gh �Q���Q@)0n QW�5w�a��g�(�	�n���sW�'N4�.�A�	�4�R�w� 0��8ه����ĜU太r�:R���w��Y��S���_�����h����o�'�}5M�AT�r$!��SI���W�w_�T�zDR��t|��)�`���g*���Y���A�!<m���I�kj���mH��/`-D|���y�q����Ž�v� �{��ɖ*t��I��H�������C�_�n>�`��Fr��l�A�����/�5m7
=q1C�^��D�p��ġ�$��4����a�ˑ�=�_��C�|w:�ʽP�c���niϞ,`����l�x:���I�^؀��
Ы�^ڤ9����-#��z��p���3G�T��.T�+4�|�\�W�M0}Q%V�!I�|�z��X��l � ���GڴU�$b�6�݁��&/N�w�9W���9=���A���D�J�f(�S0��`b� �W:>xO�+c�ÎM,��u	�;P�&�	���]�O��	St;d���B��A�2�����g$��8nl���̧��� 9�/���<U½�$P]M�p! ZQ'�
{�{ѥO�@����H���O�D�Ц*�>E�_%���U�$v��XM�g�!�u���ū��y����O?��/��7xѣz*G��Z:���	�؞�S�DH�~"��s�u�܊ޱ�>
F+���D("�RAp�-u;�_��K���d��O5ari#9�eYP�������ݴDAL��A��h��.[9��}�~?Z���M��8�����\	�!o����.^"N��+4�贏��}�w�0&.KF&�:�9�f�V�	��=!��؅I��{=��qB	s��#Hc�ǩ��`�������]���fT�ES�#y뱙�*����k��`����n
�ŶѥsN¸�h��d����=RP���4��&]�+B$�7��̰2�upE� ��I*�e9B{�Z��T��'>���{�(�&:X�=[�����隝_]J�8������g�ْ��~��r$ą2�>�av����v�Sv8�A��~V�\x���A��dp���J�r��������P6/>w���)�q��zn�kOa#�ni$n�g�-���M���?RWY0�(V��� 7±O'�3�?��؝�ݿ!ko$�n��9�ŉ�b�Z����E�����N��l�	�7����)<:�'��2@t;je�������������d��$V��D�Tep>���}�Uc��Dn}\�z�A3޶��ۇ��.���Cp�r�^g�:�U���|R*R�a�Q�yi?*�D~u���A�g@�*�cq��A�70]�I��Y���cF�VQ_{�*~����0dJ#����5o� �6'��,�3o"��z�`������ތ����E�gzn���f�*�T|V����$�y;E�k>NPpJ�R,gu���jp�Ǡ^�� �ڂ�^�Eި���
���ڗ�{ѡz?BïL�_�ѡG�I�Y�%��0��v���5�T ��eJ�h�5�'��}�vE�.i#9-����.Mlr��U���:����xE��`SSW�>�k��#y\��
C<��w���9�Zz�=��i6�Ʌ������ �!݉���U5�W.L�/I\fx�Iϼ�X��#ޢv�0K����N*;T�r~�O=���N}]�hU�)>p�+�ҍ��7i6�c�3��:3͞�TK`���E�%��H�ç��]�e
sF�-~��45\�� ���!����!�򗴡s�j��)J�z�W}D�#����@�����߻�*����%���b�1;R4�L/�xSiO��`� �ī9���n��(���v��D��k[[Ys�1sd����a�I��������L�wM�Ж<L/�Q��[4O -�?�m�,eX� �U`���5��OUr�[>�ML�tC�B�^{t�F\��\�xT"v��Ŗ��|В�StƤ��w�i�*@;�Ӳ㡗n��l:���u�n�����?���̴�d���2��-��g�-#���H�?a�{�K1ބ^'���'�֛�+A(@,�epx����4�d*�]k�h7�T8������s���X���P�i��r�f�_�Tz���\K˓��}͸�3g߁1#"*d,
���(� �Pѩ<|���
� n8<��P�&�e�p�T�;�����)���t3��^)��(���o��L���� �Mb�9�0"�d��e�_�*8�����E��v����?�`p��f'�q�A�Z�Б��j����
�X���㍆�sg�''X}1i,�<���q�R�>�0�Q��^��=ۿT�����K����Pk�w�)6A��\o ��.`�JFg�ʶ�swW�ɗ�7!��Ԫɘhk��FQȷ����+�����ү�h�����:82�S���'��|A�;B�^��oX%tN�Qd�M�� hEg��cΆX�7s�J2�dF�������8�s;�롢�uqo����DD�w>ے�ϒ{]��Ҏ�v��Og6�t	���:n�٨�f��/���qt�fĠ6��҉�ј��4�?�/fne���˳!�)h���K��v��C�*_�s�c�M=�#���Ҧ�����;G��t(ȑ�9W�ȞI���'˷!8��i��������N�匐��
o��Wv�l�K u�툯�F#Z�[�)������~���nbY����=��g�7�P%�W�1�x�Bw��I�n�XdM�e��Twe+�q!6�
�|��� ���|QW	����e�{��)P�o��@��GARD׭���D�Sf�޺�4S��WC�*j_	eᕀ�6Q7֤���+�H���K� C��G�_\-�1Ǐ\d�n�j� E<�N7q1��֛�`��~=�6�i���JRӍv�b7��I�o����*d��E$m�"�7�b�L�~�⠜}��,6 |�[-X_���,-�ot�]f�;U��3ōVV��%�PK�2,�vH`�3���^K��s=�m!��r! f~�ȢS؜�������eP��Mց\d�4��p�{�֌� §��^��S�{3<�1�����c ����0+"��D܂����!�1��,1Ҡ�� 4�`F�{���,j�H����a\�^����L�����XF������Z����������#����w���9M.Rarb�k
F�OSR��L���;Bk�D���/;*��Kd��B�O1m��$\*�50�^+y�T��yN�V!*���_nΒ�abl,��!�x�9�����l�^ z��X�޴���R���E2�V*Y����4�S��YsO��{����zˬi�<��|���a���e�=�xXb�4���	��F+\��s�8���-_F!���0�d<]�]Y��R=b�PH���#vm�N,������)���;�(?a��+0`/�*�0�"\��9]�4~t�,�r|���C]O$�xB8N��g1ϡ�����MՍy��$1趾
��Z[���Ճ�l��}�����H��$�U����ң�4�<��N���D�8�rP����K��$�i��c	�#ؾ
6���^Z����Z%��Ȼ����.�a ��
�����4U�y���$�3g��[��T��}����_��W\�?�YW�;qA ���Z�t��[�|��ٝ/f�A\���pt�qw>�o�g&C���u���f���ehq���Mg�g3�oU��?�!��yk�����M�|o�#�P����*�>1�>.�:q:j]��8��sA�쨞+�]9D�Yz�5�s���ma��۶�liibZ2��ULR�|QP��o8�c����<����
+c���煎3�sIR)9C�VEH���� 3��Q�w��K��22��[׊b��������G�d�&~���x)���r�7�j�(�J������Y�*G�����6��[]��2�`r�G���l��8�>�R�������j�
N/��$��Ѕ�������ؚ�NKaN�P��@'J�	r�|���-@��gmX�~ǳ�@��H�c8y��Vm���
�fH4�+�P��wo�cKRס�g�i���`&+��3ٛ����'��12=�"�O�Hˢ!���/�؇y�ʨ©�� �<E�6���/-k�Q�8�ҳ���a��a'��tlv�����=sz�q�џ�Ă@&3�=�����:�띁=c(�����{��l� �Zj�ɲd�����Z�QԊe�z�W�q�����`����t�D�J�`}����p��c�%Gˌ��:2�R\�%�.s��ʨ�&ѧ������Ob$����]x�m�17Тw<1w�*���U�N|~7�٪]��#����+�X��9Mg.��?י_q�;mNr�U���geV/��M�6�ǜ�\����� ��$�3s�3��>�a��(�h��?�d5����֋��s̤�b@V��bko��Q�˟�WkW[����"��o�^_-H�n������$r�`����B��LِBȏW���Z�2�"����W�
4ո�J�D������=�d[��u_Ռ�\?��;t���D&t��D��z�5W�V���`5:B�+�B�o�d$�Ͽg��Fݽ���܋لiU�~����z?I�F��[Qd�.�UF��Q���	�A����OL�I~D���LHE��7E?uQl�RV�?K.�	>�%�#�-�YI0��6��p�EU�K�1\�y��=�2̠���~+o&M48[��}��G��f^��@e�q���}�)�|Q���oQ%w�=U�ԁ�{-��b�������:�����]A�(�
�9â�� /��Uu��.�53��7���j�hڡA�Ԉ�s���h�Z����	T�F��{So�A�*+�EW!(�ٍ>}���$#����0�(Г� <��r"���Gמb:AcB���02l���x�S�N!1�f�=��T��k�C{.�-�OB��"���O1������Y)�Mqc��F��+.��s�@�u3�h6ɾ�}h�0�b�kAj��)��8�� �o�D��C:�3-��9W�h3=��Џ��Z�b�j��2�j*G���!Ae4:+��"��5�J�n8��@�a��U�*³=���61��=�}��h�W+����`V�d)a
,ц��L��`�7'�,��Y0��jy`|Oeh�L�T�x�	�n�(&ł&��uQ7��k�3zQp� _�N\&a4-|�&}�IBC=H���
wTo�ϭ�u��(k�΅���r�"��8��i&��a?�a�c�T�̈4��(�(fv[T��
{Xv��@��Xm�'ZV���J	�i�F�g��ˤ�{���C��Ƹ��2 	�I���fb�
9
5�Hh;�ŶƢBloYQE�_h�(�&��˥C�&�E��O
t��ۀ��hke_�|�'e�fυ:N٥vg��%�ST���>Ff�91�oH�]I�i$�{$�cCU=�|3e X-�`��(F�\��%�+��7B�궑� )\a�.,���tbm���S��\�Z���v`��q�)���{\�ůߥ֘�Msյ��h@�v7c�E$U�TJl�&�tz-ht-F�T(8MC���N����::�U@�M[#���F	�4<^U�tn�b�����)�L���������Y}Q`����Uk�w0n��P6�5�^04������i��ߏ��61�Iؓ�`��&�����+�V:J���\��@��bd��v@D�����}�/����~��'�UH�!u5��/|�\�q�a���<�	2$���M$q؁��jX�4�an���|�%�]��P�i�@�}�zg�����T;,�_��[%��W�x��2c�ȵ,�!�m��no���^�+ʩ`��'M�i�����F�m1t}��_5�3��+Yi4̓���-eO
�ß�!�<ia;�>�t�iȟ�޸s��Bu�/�¹�dwr�s��"U��X*9�~D�.���߻��.���?�cK]2&��꩞�iZ	T��l����Nf�^�C#�2�^�]q���K���f\}�p@t�C6�@�xGz����C*)z�������X@S���
�%������=b8ߕ���1˜d�oZ��z#x�åS�h��2���i}�@��x�c�ث�.2�Lx|p����Bq�s;���r4���rh���{=���SUt"���������!����=hW�π�p���
��q\E
��؊�y-�?LT(NIp����_�j�=V�	��8�Ja?���u�^��J K_&����%uFΛ��/~�͊�a�񵩓�T����6wb�ҩA{I���c#tt��L�Z,o�����Q����ޤ�m5�A�������2i�&�:����U���t�,.u���Y�C�(��,�ߘ8D���Y����"���ԕ���ٕԇp
!�"w\�b6���<˳���(������/�=2K�S����_���Z-��Ȉ}�I��g �r�����"NR9N#�"�K�=�C�����c�$��;��5Uh#��=��k�,w��%�(A���$����
(�c���2�s��T��7k�"��a>n�;��"}bW�K-���Z����\�e��g�s�lK����t��ab��>��AK�̅������UY��t��Ѧ8��T�؞8��.���.��,�?��b��b�K��J\�,����p��z��bč�4��zckvjF���s��Fr*��������g��@������^ƕ��Zߧk��|�T��g�'���2���_���ؘ��,�&�5���N �N;�Hq��-���F��#
��/}���n<�c�˷4,�Y�M�,%H|mDTG����v4|zUckm�b!F�Gpdv:}����!�5dMY�h�|�c�d�g�lH�x:gU<?(Bn�WGUa����_u�(+Ѻ_Z����@S:��4��RzX)��!�(.Y�Z<�vC��H��P �A-Q��@ۧ*P]?�?����i&���v���5�>�g��f	(v<�QN.)L���h5'�`ya0
J4}��)"����.B���:�v ��/�,�Y�g���B�b�F/cn|e�n�]�����z���-�1J�4o4�\��i7?.5�\ܺ�uP��dC�o_�C�V�d7Q�X��	���k�L�����{��:8���:����[)�-��;��:X��+D!s
��eB�l�
�:)���M��-?��R�B��Aͧ�&.�R���5�l޴��RC�U6 �
&ƳT�x�oJ�����L�	�I�y�5���]���nF�����2u�����J��f.?2�<�"��q���n�Ȑ$-2� Na�63B��o�QG�%��Z��!m�&�ɓ�!|ܬ��?a�1\�oh�`%�e��Z���y@���Q���5ܘsG�B5�`ɪW1�cjK��:"�;yj���X"v%k�w+��F��9�|�������{���O�3\!�6X��\)����F2�PC1���-�����`��������+G��� ����9SGoۘ�X������{Gu��v�ܛI�&d_�L.|̅�W@����qf��9�=Kؙ�A��꽺ɞ������z���ҳ;�m��<�{�2����G/�Qa��8W������2�I�L�?o������5+)��������;�Dr���6���\̽Dc#1�C[p�^
l���K���֟%@�,Nޙ����Ugǫ��esW.Ț	�	|#�߉�z��(��p��:w���X@d�L��hq�MbW��.ZD�����h=���:0�%l)�_yi����j�Jг	ޔ�O_��Cs���M������&��������&����i��Ќ5���(�~E��l�c>�/�����n2��������2��C�K������	�r�I�o?и83[��u)<��i�-�K�=��f��4zK�֍x�W'�R7CVN	P�Lp��mC�ep=+��/e�w6��ZIz����BҶ��[(4�)���̚t&���xQ,���a(P6��
�vS'��.3r�$f���U��Y� ��O�zr�yo�Kq$v'�T��6��.�t.��P�-iX݄�.��{7��34�zf�`�;�����y�zE�U��-n�Y�FRM�RS�7���+���V�TG�$��8��F��!��@�2>bdҁ���L�1�4� h�G3�A����8�+���yH��-!�P�(z��e�:��Ł�}��,�.fw�����ZvAh��TO�1�Ȭ�����m1T���d ��<��u�}� n�T��|Z�? �]�T�ab�t�EG&Yl��#=l���Һw�O\[�P�D-�Y��Cc�*_`}�&5^ڃ2t֝����	׊>��-{='7�Z���i���Lt��($A=��?̻U|tiUF,�{�$L�>8����K>�5������fP5���1��P�'���+_��c�w9��׋S�O�1?8#[�i[���^U�jSl����e{oIaͷ�Ȩi4��Y}3�9�M���ȸ�(�����Zkg|�P���	g�t{�x����-P"7�ЈM(�Z�E��E�b��I"z��D(.Xm�l�.�ﺛF@K�!��c��vU{xJ���7,#D�JJ�4��ɧ[�9-
3Жˬ^6b��G����~���OfD�F�Q�e�<�	2��L�y"���i�̭t�)�D���ȣ�y��p(n��O#J���HΜ�U���f��4��x� {������,<�˚�CJ	rO�F���Mz+H��3bW+�OyeP�z0]e��1��'���9?��.S��*A짙��l]���"�1�Ĥ/�����d�(�]�m�d���#T���pX� ��k�Ǹ�2H�*-��<� �N@��>�2oy��I�;-�Y�}�u��e��c6D�q����0���hB���_�b���/_�4�0�J��A=*^�I���X�"A�_�Zr��5�1����;��5�-VI��^K�����Y���֤��~{,�̱X���a�hd0��@��P�J˜ĥ�W�I��ݞ����e���S�b�(�, �G�\P����G�%쵕  ���*+�^Xrx��Y�&���2�p�l�&$;�F��K_[e,���/����G@��}���Wp�;��x\/so��~QB�3FxpyQ��!��"�?($��}��wr�}�����C/Kd*��
?�$$!x�]eh]�{w�吴�c/2Ҋ8bC �!ջ�QyB�|�*��"���HRY$���Y�I� ���}K�tU��4��QB4����5&Y{H��.!kc�R舎j��T1Q��s]?EF	X���������VFF�Q��b�wL�8"���S&:�(��nC�s��W���5!�T�t�.S��p^�5L�9>�<�Q{U��s�Q�7S��JnF%vb�t���17����#�H�G 6d���|�I�N�q
`)ˌ/�V} ��X�8 `�x���|u�Ej�l�;w��:�H�	XQ���q8�
�P:����.I�n� ׵&��~�z�S��R'W��ǹc�YP��|?�(0?�W�폼�9�#bfJ�o&0�@ew+1|˥���
�����C�&�
ܜ���SW�|r��Ϳo��vߝ~�����=B�2tvؿ|r���(�V,<.CJU )R������3 =\1�Ď�Wٲ����V���=�I����6W�^�w��1Ǚ(���I��*|�"��x�?���~bٴ���f�LB������N�4-���о�vؼ�@��@�|#�92�ysL���J��y�y����H�t�Y�F��.�;H-�_��g<��1��$~��_������c�5�+� �����&c��re�*&s�|��ϭ-X���.��H�ׇ�����&�:32p{�K�i�?�*�?�lLx��#Ǻ:���WG����=�7�#���G����B�b�:\N�m-�x▞ͫ@���G��g�L]�>���h��R�9����$��U4���.��D-g��<��p�E �W�� �Ϛ����7��'�>k���}�+O,�'����Mq^�;�gE:���P���)m[��6��1�a�q��Of�e�-�y>�B�%�<�8�Oi3�X;s�183O��U���h�=��k��#�W�s2�y1�8���;[m$O*GUǮ��R��)�^�`�(�B��-��%��kG�C��"�J-qf�U��-v�%�W?1ڶx�ƿ���'xel�W����u1/2��9�u1�(�E^SP7�j��b�&c��t�*|���(G�^��9(E2���TC!��Xu�Gؠ�}��_#1ֆdl���%U\�;�w0��G�w${���	0"gu[;	��	3{F������z�՜eA�:hV�}��j'��N��snu�n|r�2}� 6�go��_�p�Na�,�5m ���6b�]�yF��аp	8,.�6���0R��J�$��ܨ�E�3b�'����7�+�������3zwv��Yg�0͍h^���
�ϩI�k�n��S�ߣa�x:>�Z
G\@ ����7�/�{��.��_�x���O��'�����تkw`���0��:!7����YwX;):đ��C0X����ⲻ�sg�%�F�J����?J���ELp����68G��M7��
v��*�T���F��?Uk��ϳC��H���aw<}-Ⱥr�k�X��)��rr�q�R|!��:��a��R�Q �ܘ=� ��E�D���6F�a|�
�x�\L��<�l?v��Xr�o^O䚐<C�x�8�V.<#�͙k�a)h4�������������q�}Q�DKF `��%AW�*Z�L����rv
���A�͉�E@}=F���ޮ��s�Y$�H��������.����Ҋ}&v �`W��'�Bd3	�Ń�?��{Ѽa1���Hx�:ā fLb$ƾhB�E��o�];62�/��q�9�`���OU���1�n�q"���ȭ��y0�,!Z�y� 0l$S��ܙsX����s7;h��A?�nz�A���O7�l��
�"�D==���'zT�,��ԇRP���3δ3�j�w���Wg0�$��������;�AU����;d
t�+~��	���̝�&A��*���1�ȩ�s6.|$�Y`ݸK�(�0+GD���I�ݙwC�;�J^�����/�xC��2�5Wzl��xΦ��E���k�5��}�mt.�B�x;�����yK�I�@�J�	YӋh�F�@�\��p���1J��+6+?&@�Q�gV� ���A�Z��M1Q�Dy�җV1{BZ�X���p.��F�J�y6�L��s[ӈ]pG�qh����T�_���)�7���h�f#|�"F��H+�*�]�<l.��
��׳��ǮTm"k�"?"�8�U�� jJa��jF}������P�-�Mִ�����ɗЇ��j�x�*8@����H^���x@��x'���!���9���A�NPe~���Q��y ng��e2�,��M+b��:����^�8�GB?�ض�6j����{Qo0���ם(�5�yɘ.�9���"!e��~��p�g�}���
&H�.���kF���t��@��{�}]��k��R��ƛ;���ӤK@�'�������
���0���dO���&��*>÷[�c-��p%������wnrq�#�i��<3Fe���g��)��!�����U�R��xy�b5��Wɟ#��ː�j���R�Wf��]� �"���DA�Vk�����+0�gcw,FD�h��S�I]�G�I9`��H�Yu�wc��p��[»�Q�+����
#x�����*�Z��G���m��r}]����;�[�,NB�)DP�:g,�]m8f��ONE�I<���f��"�P�]R�a�UǏ����&��1H�~�G%;?�Q�p\�OJ�E�Q������hb��ѣ�qh�1��-�&RϿ٭�N!��=���J]�3��#Y����;1UNM���B&qiZ� 1�w�	7G��W�{�a�]�s�x�RN1��3-N���N���$5�D/uB n���0��+)�>���g�C�M�l[������� ��F�#�H(^�Ns��}����O���1�yϊ
.�+."T?2��}�&����N����[���Y��? ��Y3AɉZ�_	錣��%�[G�I��i��F�H)e�l�֮��F�n��a`�/�~����Y�V�v"���qu�+@��d>�x���{Y��m�r�p����?�
�������0>ǣs-�;ZзZF����1�f��N��5w�ڐ��`��p�3�׽+�x��{�4���!�(���j9�[sɰ4t۬	W�P�Upr��`i#@�1�m�G�?-?a�ƞ���쯄�9Oy�:xP:�ft�$�tJi]�2�6�����m�FW@Ԝ����_��2z��)��I����\�~��wVֈ-�c��W,{���Ov���2EfS���$z�����f~Y������Hߑs��~7��5���Jx���㏡4ه���~nώ�<KZOc�k�%41(�;�I�*B&�Wδ��y��%�o<c��P��:S������@�G�:z��"�r쓞P9hT{��N���CR�a�Df�{�3�8ԛ#��B��}��C ��Rb�����j λ�o+F+R�z���lX�n��A�X�l�ý�L%�
-��PH����/�|�yՃ�$�n+�h�Ҏ	Oa�
Hf6uZM��k�W�2�l��!�YM��`������Iu�?���U��lH�:��E&i١�3����l����^y ��=�g�c	`���G� �CJ�@������fe;J+��5z|Y����|�;
��L)L����%B��&�X/i�Z�j�X�hs�A�$=s�&��:�C��8_*q��#���&��d_ O�?�ě|�vxK��l�7��#��y�2!�gR�W1�4�3o�W?sXH�����-H���dJ���nt��v�RJq��{@��KT�~�<�.>��O����>( Z����$4�wB��NZ��K�@�6����x�KcE�"Q���Y�Ǽ��J��%wTG
�DR'�6z������z����b�qY��� �73�HT}HqN�*ֻ��df&:]�}�h�[#<R���.���J�*'%�>�
@\��p�F1���;�*�J��|�*���tй���gi����;K�z�!ڇ,�[�;:ӊ�C��#Pa�$mx�mb��S�!U1��,���'0���r�Mr$���z��!)����"�FY��X��6�a픀��]w�ch�����4�.�Fj�(��Т�����/3L(��~<ӹ���4�?��Δ���}_��w�
������:�3������2�����Q���1=��S���q�&�YXz�q���p�,1�-6E�G9Z���信��ZE$�N�� Mër�R$�3Bt=�	J�u��=� ;��{��^B򭻄���l�~ܩr8q�w ��	Xa��Ი�ܱd���wȤn�.WM|����kɪ0Dś�H#�����R����g@�j�Ե�_R�N�Ly�CA*�産��B��Xh2��uVQ����LBk��ɬ��kz�Y��MXX�c\�����a��bh��q%�N�ݠ�+���%��&5�7�����|G�ٛ#-#�R��}j�'E� ����`���f}'���J��WB�~��$)X��f�E�
�6�����Z⑸?�he���g�=�\������^�[�u��Jg��y��A�?"k8�r1S�.%:�Z�R���E���.��bt�t�!�v�|�}�?��/�cEJ4-yB�������N-S�ˑ0����lCzgz��{Z!�P�[i�r>%�'�6���3� R�Ԙ<�.����.��|W���74���C"(�4���v�'YI�¦��W���i���^�dx���F��`3�Ă_����}�`O0�H
Th:Ƅ0�bȵU�yR p����K����=@�Q$\zS�Gi�XR�5��H�C~��i��kY�#>vF2guБ��>���y�m,�b���������Y�C�@��D'��`����Z�I�c��Q(+��P���U>��3--��鵉A���"n�8]�|�Q����Φ�n;f/.�tJ���ꅠ��n�h�(�݄�N�ϕ�ʕ���0�e��t5���z%�Z�/|���n��m��ni4Ƥъ2ɂ��i�Β�����D����g�qF���2�<�Q���|�<����$�ej�P�� �C��z�?�ĕ���V_�ƕ�%a�a�; 7�m�v�)��kE��q���č��[}�s��H�A�tB
�u����9]L袥*x)$���R�3!�*�_$�� k�2.%q)��͂x�GDh݁���v�q6��a>�rw���E����h�=M��g/b��X�ə]�(4��D���8���8N�d��Q�@�J�Sc�@��s]�e��)�s���ku�I|3���a\��`h[�m1!�"0ƍ&E��C�OfĻ;`>�kZ�Y���͂HY�HP����2�"���<XddB&z"�|z �|֗��9�]c��0��cBѕ�b@�F�a�{���	���������^��d#���c���(�AVL��&���9ė���bX����ƤY;�]�}׺��}ӳ6��B��w��̍ _����Pɟ��d�|E�����5h/���N��Hv� �<��Ǥ̜�y.����f^���KODZ<����,�W��Hߦa�Lc邪Q�L��kz��ǯ�A�8�	��x{�!��T�X@ BHMV4*��"�ݢ��+`�����ro�B��sY"�'�>�$�%h\���Üa�1�9�쓣��p���vD녃��j����=c2�	�ǩ���<���,2
6͗��Q��ϱ%��|�ld��kW{��D�{�@ԥ?���P`��3��
>V0wlWu�*�8�(�8�;
) ή�(��e��z�vHggq��B���39l	F�w.4�e�t{�Ƒ���^�sl��t$�Hg1�*�.��)ZCY���9���'ɒ;���/��U���<^l5��d�� ���������s�0��l׏���5�O
3�!����������m�S�l���Bh��#���̮�X�#���ʫ������(n��+O���P�=ü����@ٖ���ޙx[�N<�C���A�O�T��#ᩣO�Xr3�	���h`0�Ǒg<y�#�g�Ajoo���I��	��6�.�{�v���8��+����;];��&�z�ɑ�N\�ij�`�^R��>xV��&�r�݀��k�Y�iK������)�>L�O�;�^�&�Yg3�䭫R�얣f�`)T�4N2i�R���#���R;{V�cc��&����ߓ/���_B��$�3�� # ��W�D��i���Ӗ��t��2s�_��5r$D���	ش�ȴmLD �l[I��y;��o=�!�
��<q�@/1Y�+M��v׷�3{�`)��i���5�^���2%��@�B��	[����c3���1eY�l�^y\��Pp��&�+�#��!3��4mH��ge����(-��b���U�nԅyl�=�*�`"UK��q Ctj��nz�,��=�./���>ܜY����HJ�^5�iC��b9mK0��$�7��x�G�K���L^������J�ظhR[
��M�op�m�IAL��B���%�W]����s�ZRR��H�>��9�hr꼮�9�I�	�%�}�Е
'����9�^������ٷz2�'��c�Z����9�ysl��TY�0��*ev�@��������-B�}�n�s������� r��q�G�ŗ VG��:�u�S�J��>v���Sa�#�9�G��lr��k�*���Ĩ�*j��B��I~;6�P��X$6m7�����]�_�Խ	��P�?1���v�2�Ѩ֧����'���� 5��5gWr���r��m�E3"N_��R9�$$eL��Po�f��� �-A���i�·�}q���M�R=�m��C�*��.�����-�M��r�.C���>^���M�.܌:�Eq����Q�_�E���/29�ev��║2�ƪАo�� I�"b�0�m̚k�L�b�gu��ʥ?� E���ޤ;|���ҩ��g��S�
9��\�i"��F���N��F�6�m�;	�r���.%��1��������s��m2�3�6�v�	륪ݿ��&DF*�@Jxx�Z���)�-C�����sKG�⤲D��Ԙscɏ����7��c��A�qɲ|iD	FwTQ��A9t�Z[�E�F������6v��x��d�Np�z���K�������H} �+��&Ĕ��	)�ڀ �b5�j���pQO\��Y��� W��L÷�vx [�}e���(��'.(c�j�����=ԅ ��:dc��x��V�q=ê�<�ҚZs���b���-�y�M�߿�N.�2���A"8�Yh e�J��}�$b_ݰxh���ڔ/R'��$�:J{㩂�=�dB-��s[�@�J�Z�Z�5	�qRVsV�y��^��Ȼ8I��
J.#"��UD���s��7���]�
���h���p��y�7.?5�l��lROi�U��Y6��~�L���w��h���<��,�޾&U����q�ʖq$g`�3�>��m��e��t�lF�s��{p��U�7�(׈�imjs�/���J�Xf��f��;��f��M��@p,"w;�v����y�����o�
J��(�.� ����`/�<R�:Is�J.��`D?T�lK�k�3ڵM;��-�=�~��u������L���5����f����{�q�|)�0��w��Z���݄��AX�����1�5�bo;8M�ec�����sd�<�ORV:�2M.�[��~x���˚fˬy�0,��+Ք�$��m��=w�idP�O��Bm���iea�ۙ�)�F��7�	�$�S�q�:��يE	dR?�GО�E�/yNW\9Z]VR�/_�5�|�Ц�pV]��I��wY��E N�!�ތ
 �m�����J9jM~��J`4)��X&����*��Q�����kR7�!��Iⴆ�w��6Ƥ���3�L���p��u������MG:�����+;ڊ[��>��ԳJr��.���������ZBN�
P�9�t7����1;y�L�yQڴ�'���"�Ļ�!�zp��ļq'�T��	
K����	z}[Ŗ&&�8� Cw!�~�|�{Ή��TōB�35�wM.-��#��VU۟��zm�H�G�t�� �d��T �f9� �|qHD}P	~{�������h�d|���v���d��-4�8$��7b�Rjv&���6�5y�TuR�|dx:-^,МGZ�{��-ޘBZ*i֜p�tON�g�	S��&�>0�N�w���r=e���.P�I( )�9)�{�I/��*�,L��0�[�ǀSt?`����'y_'�.L�d�F3M���t��0R*��뛾Q$��s�Փ�Y�����Z�C߰W\��FcBk��8"�m�s��B>��X�ю� aM�d&���yI��^���+ǧ$���n������|"�P��:�ldL�-`�)��	�W}��9}ȸbz�3���Ogт�쫶9��"0���kr$
x����H��N��F.�!V�yn#^輖�Q���CVO7}£��d�3u�f�q��Ł�tp�gCK��?�~�a{}(����l��:���_�$.�v��j�8����n�����ЅrY�Q=�o1X�-hzO��M���I���AU��4��nR�˛*]&A�13���F^^����g�7��H
ی�z$�M=��I Z���N}Q'�V$�N ����J��� ��~���o�����3[5v��Q1R)ByUqb�i��T��i&{����p�~K�4�,1���Ĝ�.��2�Ek�M6t��t�rȷ9dw��@ ��86Q�H����92�ƀ��	��r^+��+��+�:�b����y 1Ԗ�Ē�_2��)�O��FPA�6�c�%<�m��۽�J�����;}�2P��V�YLs��՚c �8�OM��{[������؝�=+�4|�9�����^hjIb��=P����Y4��b��2��ߨ�k?e]��d@��k�U�o�eM�<��b���3z�|T�� �)�ds��J�6	�\��~ԁ�Ӑ�^#O;׾I��8'����5V��ޔ!�*�U��Ŝ���B?�imuNn��*͟�)g��O�+�M�ж��<�#+ﰲ�ˈ��d��8l{0�!=����'�L�%�`3����m?�� ���EK
5�?�Z�UD�\o�9��1�������d��a��W�tS�#<`^�#"-"�x:� y��9��N~+\f��9߽]�b�������u1���ˎcl��x��bm�U[C��s����ߝ�~���AC�a-��Be�����$�=�ڣ�uv˖H-Y�AH�C�7��?���6U�ł��ÅS�:э�".���A�L;��6ץ5m�B}'S�QmŏG$��<�a\����8��	|���֘�|q�yx��#��P!a�Ֆ���)Ep~w�,
$|�������g�I���5p!�>��D�mM����%�J&��VG<���6���Ӕ�3�lK�i�.gM���c����CQ�>�y(��}�C]{�tؑ��X����o�ե��A�d+Y|NYv=����q�K�A�8�g�E��dh����T�V+E�J��*.Mr>"=�/ �D�\hW��l��w;�\�%�d�Ҩ�V[��w�dS�����63��[��z�m�v�F�����H�tU�|��wo2{	��G�Ǧx�A'.IԽn'�qRKH*a9�=*�>H���&�ux�?�߅� �1�P�e<c2�L��%��y��t�@���I��2n�{.�vێ�B���k�V�r(P(��?��B����;�;?n��dr%�0���f�t�ɳTq	�
~���q�0K�k�B@�H��-�����+��eKPQh� �}e<0M{wak��3��>QS�q0���|�/�'�3P��o����T]"(����8�|֌�P�	U��|(%w[�i|J4��R'`��?ܤ<y�č���_ʍ����ci��i_'	�����i}~�n�+��M�~0������r#�$�xHo��Z�ځ=����VX���ō���~�6�W���t_��O��匍@Oi�c���S��EB�#
��^�cR{Cku|�*
�0��K�Z�����yc"�901'���!�)R,"'����Q�Q�{<�4��:�|̣����B�m억��r�GG�ڦr�{|��p#����i9��v�_�����}z���f�g����f���~�+z�#>��S�!HV!�o4K�WXzi��H�5#_�o���A�{��jhL����Tt.�D�B�^_!a+�?�^����w����1���jE� f����}nb�Q(����2�f�̈�}	���@i<F"}V'N�sx�������o]���ȅ��:����9�Jae�(�h��ۄBR���4V?�>���l�"�ê�w\���n���Ȧq��5���(|�z�F�0�AI�)�2���҉�^g�!'$�E�֗�Hļ>���#�u5h]���=��G§��SG(���u�<�ΌgH�42�;� ��Ȅ_B<���i�&�8��	-x�o�{kn������>����[�%�#5+
�6>�����O��W�q� ���� \���}�4�D�!Vd���"lD��$/%���ϫZ�-p�
p��|������vwό��� q{16�s�������Ajg%���5���^�gJ�j��Z�a��GE����OO��'@�]gX|��߬�oq��.����ϖQ�(x���`ȼ@Ѹ�*���ތ�w4j��8�<�����3@E��E�59?��ֲm�7��7��Č�Z��ե:��rRth�_o�2�=6�{��\�Yܳ�V���:2p:(c�/���|Z�z��*;�L�5h�ď��q��?������`�!����mZ�y�6>D��ׇY��1�i,}����B7�!�4���DS���f����812^�T�ʤ/����)���f^B6��QZ�r�I�r{�(cԝ*�o��&M�/}�Lk���8�I:C9,;�9x���yR�o"}�����O����(�3z�
(I�
dy\p�"L������K��6u��B�c���!"��v����
�ca��t��-�ɜȗh�Xipi�?�F�{� +?
'��6�O�ئ�G�4��lR.ݱ��eD�d-%��ԯͦ��!h�Ƒ�׸W�;w� @ĸ����2y�����v6B�Ka�-�g{ ��O��a��p!��5����e����!��'��y�1*&,���0��Zcib���R��r��ϰ�"'x�j��n��7����Ap��
��'{�Z�d�´�=����"�$s��a9+$�,��LS��A����yn�>�Y����]�sY������Χ%ތ��+�}��PVP����}N�~�d�z��,��nu��]�2t)2����6��\d���/j��з�@��� �c�\���ۆ��ˬ��~)w8��z���@9�&��x�r���������mqт�N͑�U�h�����6���7��L��#�w7B�9(�1���14�+/�4%���$V�S��^��R�*��L1�A˰�@���idm��=�Y�j��~�o15��YS�a����6�=����-���~�a����h�]i��~¿�1Q�6L��ī�K���X�����ldMjGIU9�2ܢ�)�^R`�`,��0ת�Zݾ��az˲��4Z���B&�%�P<��E`�JH9���b�'�"���Qt��������K�M�XS(�6۳�f}N�^D��&a���H���p���|�'v�BT��H�ӭ�Z��4�`4�^�������Q[�>*�n��[�H6�v(�M�1��?���}��ٌ�'��|�ly���϶�4�g��[�)�R�
������ي?(�~���W|��d��@��ěk���c�2m�v"oΈ�5#:y����Zx'k�?r��8�^�W�BX�>$��b�����v
�i�dDKB�fշL-é`EO��z�4�_����&/MO���I}��-,�!\���Š�����D�����g��U���kÌ.Q:2��4m�GX�����߉�º��
��^7|J������	�#�COR
=�B���!�75���]��%KY�p�E/^nX'H�t����r&�C�rߗ�:ל͈��y7��њK��/,���W}\� !�ɷ�?�t��n�7���=��j$	7��w!�+/w�byc��5��lDka҈������̅Ǡݔ� �[3�4D�c�~��� ���Pw5%N_����_8���=���?�t�"N�hӸ2�S2�r*b7��4߅��H��t�"�����fq�MN���X�F�W��Z??�DQ�@NR;LZg�/ED�s�O��ʸk9qq�I���e]*�H�.�1:�Fa�/yǞ�oy�)Aj:�H�Ws��;�^��
N���1�"YS�
)��6���$,&�b�j18*�v�T��v��8rfs��x�gri=H�y5(穔��.�萀�8Rra�dY�|"��e�:b=��O���s(�o�/w6u%�d+�i'�̷�;��;M2�菠�,o��w)}���m���i�":��yC����jPa����θj8e��\��,�v��nIkt�3t@�7x�"�w�5 {���;d��� 2b��k���?@�Xk�����Q��!���1��0�D�4��< ��#�8�f�1;Hv���.�_7��V�B���]ؑ)�-X����'I�hM=R��`c��rfP�(a?k�D���N6N~MI�/���+DM��ئ�dupo}��oa����}ch$��u��i�ylpV���)�����㷙3��B�kw��/��qL���0[�&V[�	R��<R���cf1Y$w�P6<�_�bBZCk�F0�6���!W��:-��|� ���S�n�ç<�0ݸ����Q%�k����L�.0�P�R�	{C�r��E�=(��f�� ���PPY"qQY9�4��7S��}~u��#j?����\N�u�9XnH.����'���W1��y���g�.<�Vu��J����P᭎!"A��/s�=N����t�tel�.Rλ�:��ʰ����Y���+36[o�c���R����"���8�QO#S᧩���֙�V�d��Ӱ�6ݪ]���[�m\D����@d����0=��N1��T�i�Ӹ.�U[�CP:f���>��Ѿ�Ѫ��N����h��
��|�:e)-���lI���|���XZP��b�y�;8��Hp���(�L�-������?d?;�FV{Cg���t7 a���iL��2�����&����+G>�"g6�Z6Eq%Ot���˱EZ�&���4�gd�r@IUL:�6�P�$7D�
x��<'%�R�e�[�"ɺ_��w�Wwf�h Ò�`�>��e��J���GeԬA�Ĥ�[\]��e[�UZ	��i�d�P�p�Ԩ8�	8�5K�J@�_�j1�LI�Ub?��x���8A��+\���$���z�������,�]+��@h��вA�w�$Rk�P[�^�Ԙ�4��bB�n `מ������_�p���~y���k�fF��s���7��G<�΀i襣���,�9�Kf�1���8\�!^��[6S1�:�|3�x[�@c��/�=�)(�IwQ�=�V��CL6g]��%�i�h��	�6t_P�@��ł7��%�|<��3��:�-dh��z��l�;���-ձ�Na��G[�pK0�5o�*��(��_��UN$=z�QǠ��a��2�;��3�UA`[�N7���B|d�8�S��4�W�^���%~[SQ�"t������:�3X�}���S�>f�?��������{V��Sk�++��u���o���>�֮��/X�,dN�/&$��͇�j`���+�?����́�0����:"GS����[p�B���D����<Z�����8B��0Ơ,Cp	!k�;r!Oԃ:��F����OoUY�6;�5�իn�n��p�/a����1b�DhYD����m6�K�BF��� ��]$�7@�
Z�$h�Bj�/�[�n�C/kO<��&ںBBEB�6�M4��'�\p����`�1;Q+v/���u󊃧��n���s�c��ۑ���)�M�F3�s<v����`I�x��8�t2qcA�&��PȎP��>����sn
�r���%�HH��=��r7w��
BM lOm���]���DӐ_���'���t}����%gl�z:��j���w�]��׍��C�+o�����eǌ��������*lZ�������sj������N�h�g�%7 �z�����
1�!��:�xUwN*�BR[M���0	�����^�E�i�Xwc ��c�\�Tr��Yq�!���d�f�?8f_���u� ����=�I��g�傽��Nȋ���F��L�?�-~����!�e]G�M�v������n���R_�1���kG �¡�!��T�_B_�{qt6���8Ѭ���1=§��.P�{�������4��B�y����������K�Y�C�,���C/,��v��י��i��~)�:5���$��+�jˁ[!h�#*�)���JԼ�/
i�Z�Ņ,޼$k��F�5+I*��������A���K�jb+&"3g(a��^�� ��nK�����:�*óIW���5��huQ�p)��L�%,��5:����%h�+	1הl|_ ����n�J��fS�>6Z��3Y�F��aq�V��
�ƕ��8r�*�oQyi5ڣ40w����rWkk&,)��q�����#_��\U�r�I��z�B�$|��E������8�&WU���7�e+U@1�c�9�︸�괰.���.|�Pvpw��fC�C�"�y��!�}AP��:�}�Ţ�0a��'�|?�K�ۘ�u=������_�Y��+Wք`3:o7d�h�a�����p:(({f��8X �w���j
p@�{=ʉ�拕�@�*�"k	�p<�!�nM|=)ò
��ԅ:�.b@�ۗo(-��L�?1�}ܙ6�s������o�x�&_0l>9����V���-`������[�W�ئ�VE�ي��튴��ʂ�}�˥xjQU�S�/�j�>^���ōhv�8��*����BB������~VImX�s+ugS�G.�V�n�8
�Vyg W�Pzj@��g&�n�←�YmX-��Nt�A{�̝�C�\��2����>�z�{iΈ�u�b��e{��*k) k	�r�\�J����7G�R �"^�Ghm��BA�W8�JU:�ӹI�Z�Y���T��s�@�Eʲ�3o�	�~˗IJRѝ��5R�H��ߑU��̳�@�t � =��<��Y���: fO$ގ��`�{3	���ޯ��?�`�8#=���vI�>���pO<x�{��K�	�"�YCڀwl�|��*B�xvz�X�s&�]N�U�S9�`�y&M�ko7�6��Nܵ,��#+���b
W<�%9����r��E��#��y�F���i'$$�Pu�����|���k��;l�6��t+��5X�BL�v\��o�͎�����MH�>���xĄ�H0��n�����Ѭ��Ez�gR���L�B�.*e�r���d#rBL�U��_]5u�Q��c�f��tn��@�`s��i�S/^�]h�6)�zܤ�� b�����Z"6�w�B}�܊0JvyV�����dB���&|7t���
<Ga?�2�F8�e�E�J�U1��t.}�)�K�60�cVƞ[لo�H��y,Z$LGW���߳�(�R�t��� K�0"�lu��-�gx�}h���ib���{#7��F3u{�hkmO��E�&���s��\6&����� A]��o|�-P�i)�
l�ד�C��bU�$g{M�5��IΎW�=�3�U�;�6��:kmu�VHe� 
��2�����	d��u\^yEy�f�u��Fh��5g82�#�/"�c1�:�%� w��_�D*�h(e�㮷�`�uy�</u��*��d�?�$�
c�D���ԫ�=Re��d0j��yC���~ԣq(�)����7"����S�x���䐡0��^�� ��=����+������\�x!�P��iF��7���ߥ�r�֋�A'촪��	m�v��x�|��+s���ݾ�l�d3CYf�ٱܣ�������B
a�׆T��Z%2�!~J��;e-���?;Rv�w�m�T���i"����j��nzE�4Sc�Pg����ڕ0��H�{ qHF�7��B���R����(O	�hM @�ly�&Դ@����}��d�q�r�CX�L&%��X�cnH:ܴ��a�7�g��p ��w:�=�Ȫ�qnD|�q���X?r���<���"[�ҋ��G7�x1x��W���ѻ��^�T�D?�Am�t�b'"\m�v���7��W3����ki�-�]�B�1r�-)z�XM���|	��.�1�FK�K�����%S���b���d5Aˏ��F���a�(�?ZR��At]*�Ĉ0He��mjV��8�O!R��D7���ђ�Đ�bJmy<!i\��$L��]O�	��	�0$�|�zeIhz��64���_�	?p:��W��!��y0�.���ʏ/hu7���ľ�-�,x-jpc�P��#�~�p=7��(�į6�]����'��/�6s$v�c��a{ۑ����J3	\���2.;�h����j���|�b��J����1��C=�q���W�Q�SΨvTA�YO�����{cr�\�βm[�{��=\�_dvh�H[�2��$��?�����j�����ro����C5�a=񞃗�6�Qp�kY�/��e�vL�[m�3�ƫ/�,�dfH�����刍�̌h��g��5�3�i*��v�?E�i�]>�,��Mz_��

j�<�ї�i�3T��?�8`��?����	��pTm6�^m��>/���C���/7�ͼ����A��+P���,��������M��s��j�r&�Q۽ۯF��5F��\������j\�#! �Ϫ���|�!N�x�Hh��RY��ʸ�a� c�}2�m3�n@K��D$S }�Z����gd_�|a���3�������I�2ve�2�t�9�{7/<�X�i�4i&�<������~��*�����\�gw��n�g^�P���P�n�8��d��:Ň��F�#�Ι���2�\Q�j� i��`���@_�ai����,e��R����k�e���V[�>b����,�+��/���`�s!*����Ƕ=�DƏ�F`�=���_�J�����Ea�I���XXj�zߪʎ���,u~�Ѩ�?�n'��}��Z�	�|�w��m(k@�^3���5Lg�j�.^�KGνg���>�%(?��z�ِJ�e��Wu0�;�a�y��1�K��g2��g�����,t��-�Q*!n���{K�y�|W/���q)�5M����HJ�b�1�dUn듕 ��F8?�yT�ow����4+7mv�q�� ۸���먱�G�U$���<U�t�� ���8�����w���(�f���Uy� 3���[���H�ϸ���1a�!������´��l��/tA�v)�C%S�Pv��X5T��!�7"�#��QI�F�T5if$nm �k�n��c7�z襛2:A�qVer1��s�a3�0n�Y��}_���ɇt�@$q�<i�Xw��IO'sE����f��0�H'n��&�,>M�a��Q�)�-�e{��J6Z;R�xO�CA�CwZ��!�[�3��R����~�8���{�3�*��L*����B��|�QR�%��K�q��Ee��8N�j�=즹S��>�����'n f��71��h�1�i�N�lk�������j%T��d�o�C�v1�1��ÿë��HQ����.|��iHQ%961�r�~Z^��y6,r�\�)��i|���� �\O^c	��w��qt<&$H�>@�U��0^)�S;�h�;Nɫ ]�TҬ:(���F�WF�V@�������Œ���cڗ9�S��Q��(qX"u����B�(iF��poa�Z�r�C���j�Đ�{�� �O(��)�˛�z��]�\e�Ԩ-β``r�P)�x�TRTgZ*^�˦�5=&�?�!�0���т`�����o��A�	m5�+cJ�e�b��*8�)� Jh���<8�N�d`V_ݘR��^��CAu)�P\�%�c��wל!�1�x~�S2��V"�k�:g��¦�>�0t�G����"(���9��0��y�����>O��H	�!�7�ݑ��� �aB?un�),�>�K94&��Qw� Ƀ�#!s{���QW�0_p�.��L'OG� @��A���+h.米5�u(OJY<J���
�'m�ϧ��U�8N1lk� 
N�Y.����v
���Q*#l��m�
�g/�ڨq����+���������#�����3�鳾e��LN7��iUm���qT�O~[M��?$=��F��E��?Tݙ�-�_ݨ_
ձ�:
�'B�r�%3�������*��@.��v�d>+X�ǚ���2�>q`���pl[a�h[Ui�Ǧ���V�'fu�qN��a�R���M``x��]<��z�0�x�+�:l��9 EB���>f��Z1�47�|���y!r���Ķ��ѳ�wI�]�r�K]ă��_��}UAmiy9(�7��4���hV^�����r��W#{&'�Uފ��v�$$���᝘	&gg�}e�5�0���&�N�I��k�䀦4R�E5���D=!��	����E!*���$�j#��i5����D.}�@kvgė)M�x�ë��3�G�e���Wn��r�&����?�ui�q2��?�J>Gn���ʅ��B��}���1b�d�)��}��yX�*3(��%Y0��_�`����h�P�l�4E�_m#gs����k�YEW�3�7#��
�qᤢ6��(ۑ�����	�>F�qܺ��ϕj��߻��ڜ$d�S/W���"	����ŉ��߽vml�(X;?1���i�ix�Q K�]$�?��M�,��e�@,0uF�����������n!��Lw��5��. �eD��/J��Y0��̈A�:���U��I��Ԝ6�)R� V����M}w�e^(���OE�J��SgʈS(����+y�_2ҡe��}��s��)j�&�n%�d�J�j�vosR��H�d��svi<�`1u){Y�Mϻ���ّ�4W� PL¾o,e<'j&�F��m#W�'�D����ߤ)3��t��H����@۸f�u���R�d�<z���&4/�/<K�ϕՄJ�ȏ{�~�T�"F}�E�8��_w4��$H3ae!��.��.0�!�f۾����������Zs'�X
�W���݂��g)�����4ِO�j��tEq�u���Y�Dz�{�e"�Ḽ��Rة�I����@v���P��axl�;���fU�������������Oe6_O'΍��)����0�[�1�Bd��aThȖ2�k��B0�����)�vᑱ�Iu7�A���G�d��0.�Cј�}U��s�ٱ�ϡ�?c�*j����zvN��L%�e�X��֊�!n�-sUй��P�jd�~�q�i�o�v{���;1��DKєN�]�>��q�Ԫ�`�c�9q\�{iv�g����,�|�-5�kTe�ڼܪ��UB{|ޣ@�5];)\b�1�	�Kf��b6�|�bi�;`|+D變u�Hi<�r���Tn7Y�����V�ݥH�ʁrn%0mk�ӱ�ژe� �L`��D-gLƄ�P�N��R^;�#p�������{���t��r�I7� �Z 	�q�#�V$���A&k��L�<�O	�ھ��������LrWE<�=ɝ���F�eT�B��Q���p�����X���}��I�R³v%�'��94���ѻ��-�3wu0GҔ�x���~;"�A�
t��
iڙ���NW۸譻m}襮*3�e�vr��I����q!Bp6ăޛV�(("
Zy	�6Ic��Qʂ�&�e���hshc ��Q�6�N�K3���Q�����v (�}�,C딫�Wg�o��G�ĩc�� �93��yfN�1��pmZ�)0���� �[E>'2~���J����y�L�A��us"q�(�0PC�;��(0,.��dn���uJu��㔃�i#���I�Q��y^�B�,�6C�}%;́1��!�~��Sq���N��ⷸ�=kQ��;o��U���J e��Ћ _ 2ɗ�ïg�5��8�g�Ya~��rH�E��:�w�ͦs3�w�_�d��M��K �'�F��]sGy��f|���&�h���e�3��&3�gFX��4��*o�z1$r�y�VM��)�L��5F6v�@�����tÕ�������E��!�^ک�đ���Oઝ;�f�.��ٺ�!;.S�t���$�.�\Gt����$x��;��ag����0,����tnq�J�W3��@�F�hz@W��]����(�.��<}`���&Zq��47�ꧾH�u��e~�^�o�.�Õ���=��"��M�B)�9��B��R����\$�<W5e]X>1��aY%X+>THj�=Or$��H!s�o���1����a9���;;�S?p��Nrz��?m2�Ed2���'��i��A&�R�h��M�F���tPG��̂|T��oc�ۑ�@٫X�>A'�z�,��+��4P-��U?ꫩJ(���1"e�¡��'e�y���D�  �s=��0����<�x��I��N����&n� g_l�`�_sf���A�M���]{��<e.�#@a\�o���Z�OU��q�(���ʼ/�����m�?77> A��O\�w��v��'�)q������-AlcJҨ;~x��`{��<�Y�eK)|r��f�G��1��'�Q11k
�yh���7����%�)�_̐C�6&�֟u�ɢ6h�۬`*}���%� h��G��������̠xP�?���w�j75^���vQ��40i�BHG���S�^ė��l&iЁ�^���e�3�����;h��(q����:>70�oF:@ͧ�������c����n��ƶk��������t�<�YA`W�0��Ge��ty�D%�هo&�u�=�����d��Ͱ��͆���D�[�E2�ӟ�]�Z��f�B��r"������՟���{�����������z9|����לO�&kAfPV�랮�E	����5労u�y?��RomGX3�������x�b���ՓPK�!�70q��
�SH���7�^����g�,yD�C�u���2��<��~�m�PTѹTO#�'B�+[�k���Sb.6�.���ʼ�S di�n�*�1?� 	9N�aA��%�'{ˉ��h� v�������M\�Tl����4ΊS	�����i��Uo�ِ��4=
���؎"����6����s����
��x\ }a����������֞�RS�O/��s�߲簓���B��2	���i�G��)HB�i�避�R�zLz�O���G}�pbg�m��V�Q��/���A���2_cB�8
�q�9�LL�9�#hL�zh��I�~���_����A�(`z6m�V�"ح�	-]����զ�}����_P]�(�ǣIVz�ٔ1�+�Ӵv�N�X�\�x�8����gDx-m����V�Ai�s7��O$��n�6*t�w�4~�fX��g���(%̒�9½�kw����`//����ê{��a�Ѹ���8�Q8D�Ӫ\��PV�����õK��5WG�Aɕ��%��t8�.��K$'�L��N}d��aTO;1��]�S����/��J��;:��X�s�f����$}Pv�p�@�,P_T΂�	������s��o���g0��j�7�� .M�4@��7��4�k�qHF��
�MHyޒ�����9��h���M��&](��z��@�Ѫܹn�
�^4e�*T�+�;c������]�'r��\ �$��0͗P������h��H��KA���d��V0}Rpv�rlS��.�zW���p��zB�v��L�4į&��'=� '��yw�5��im�g���Oc	����:��-m�%[��y���R��B��C766eF�u��"+�w�*>�Ըj��R�V�4kdk>�"Q)ך|w����ܣ���9��Vt|WC��m�ogCA�Ĳ��5�`M�mARW
�
��H;-tS�;���^�r;R�x|�H�_~�>�`@pU�xҗ�#�0���l��'ClG����>�T�` ��	]�����o��zRA_�ISh��<��|�X�2�b��SȚnN��#�	���=j9��s�X�k�N촭^-������lܨ �ә��B��3�R`�F�G_��n������8(>{���5 ]\(�Ҹ8�2�	 �xf�	L ��Uy��=�)@&�,����*j��0�JjY��]2�+b��om����.��"��������9�&�c�!x��n)�x0���p��_U�|�]AJ�?��zSW/�å隺���JHY'��b}3������훉�5��R@rB�A.m	N��px��(e�	��嶼���3DBڣO�X���H_�<�;�4h3�~�gw&���A
�����~����x�����L�>bཞqW9�qd��*Ъ��^<ʮf[��'�z���ϻ)
G]O�Y"�oE-/~>��V��`�`�T��9UL(a�����C�1�m���t��lbWi��L3Î�͈�6i&1y���A��AQ'V>{�-h�f}E`�I�Q���I�Nc2���;8�6��a��0�#Btj<��J�gftH/r�r:@Xi�����\�;h�E$E���Cg2c�_�v�����]^��1Yf!N�4�u`�,�YZF���VBg@�ㆊw0�F�P%K��mHD������XH4�&s�k�Th�U U�ruڟ�$�m�����g�Y1���wq�_���0o-Z&��1��5�R����vв�`Qa]l�yc��`c�����S����)�
�5ؔ���ü���,~'�qi4�g�G�;�F����z����b (O�0��I����a���\�<qɀ�� �b'b�O;��o�9��+r��K<�M�<���H�T1t��-XRP�3��]q�� �Ç,�N�����ju��#T�b �j��A2_6Ցc��T��(����I٠�i؋�N�/�����_=��]E���Ѯ�c�M^��C��X0�X������vn�$��ո�]Cp�JO��7�b�}{��R���4_��q���f�34���K �R���a�LcKv���giUR�\E��f���ar�E��f�������ȤGɟ����k%xK�|7-,aW>H�e��ܞM{q�'x�uW��W��op��xll�F�nwn���������2�^9�eû�<gJp��=`�t�b�:Ս�Rfjx�@	&�7��OucV3�uj�t@'@���;�la"�L7-��� �mhT)%�����a�G*� ��Ja'Q�Q�r��6�u��r��%!Q�U���@�v�^�ِ��f��=Y�����)$Yb��%6� 
��(��r3����<�^V8O�X;���C�7�8�}:���E�p6�,J��v8��۰,��K���Ny�+pۡ[OP��{�_�������̌�7��.X�#���b˽^6�zX=T�f�ϱ�߹��!�Pu'���j�����Wτ`��&�!�&�}34���98����/;��{gqm��@��^��ͪ	_f{c�����$7�n���%�e���{�=q}�i97'Q��I��r�H�iQ�S|��^�yK�X���ɱ+M�Q»�e���+�S��)6�����<]?3�����"$�%��5��(^;����r$�M�-Pb�劰k�c�%V�6����ip8�	7�5�����L��=��,YJ�����%��׷~�0�	V�w���d��x��OA�v�8��n�z�T�E7�����G�5J˩�<��b<_[c�Ƌ�F��g}�_����i�^���g�0�ܒ6g�����g`E�	���F�S:GFr��
-e�:q!&M�Xf:Ǐ�\���]�4
���:��eR��J���4����veE����V?�jQ��Z;�oi���0L��Q����A[ �_��S��8B��(oC��	����a�s��ti~��e����L�Z�ѯt:�Y�A�!�ܳh��Y�J#\c�7��y:�p��k��wʘ�O�ZB�h�cpc(��`,}K$r�^v��*h|ud�/��Ln�ZI�MApL��Ϫ�V�s?$	~���Ə�����b� �%��W�/�$`�C����Il�W�nh!î����M4���� ��5�� /�$��"�F"3��n#��c|v��	d�7����_�=UO��E�[�ۙl	��y>��w��f|�ӡ��'�@%v�͌S�W���ϱ���fװ�|��ú��({#�~��3���؈3�0LNq���OEF�xu�A���q"xA8������{�(����.�k;Lyf�I�b����������Ʀe��ꩢ ��+*�-��K�_���|��&zN؜���$h��̚��z[�[���@��֑��.O��ض#gc���n�Y�]}�y����@/4k}&e{�����1+�^7���Sjc�:Rj_+�DfR�cۀ�&Ry���$J� i'�3#��"�ck_�߃aZ^���h��pH���szT��0���AO�����ɷqH^���j����T��
X\���@���ꕱ�Ϝ�q��R��f�C��-�˪��qέ�O(�c� -
vkN ����|^x�@Hf>'l�gu ��X�R��m��۰6дfam���G_��L� *t8 �_�M��&�������/�d&��}��O��K��4Ts�{1�`��R� ň����eE�%[��2v�¸��T�)������tj���/�j�YYSL�BqZ���w�V�,+��. 2�yx���k8��Q(�.�ͱ^����AE͟���[/p�xi��;�l�67�^s�O���B�De5��C� +O�=T���w�+��
�5H�T�iV�Ȍ���r�?!�����Yp��i��8�{Jetu�붯�ۻ�7��lgw���4�Ԩ*7m_�����0M4�^5� � g/G0���L�|���&=�᫺l���.p.���T@�!,�,����d�:�c8�z�q�=F�H�zʰ6,�(��*�͒��.��z��9��g��v�O�ٴ�lAa�VJ��@�t�����nAq��~�8�F:���B]U@�a8M���xV�.�y�ď0Y_��㈙�d����Jn�@�R�:�N_�\Ԁ�fw�}+Tx��Ը�RI�%��	t�l���xԌ�Rߞ� ;˞@{f"�ƎQ�0�r�v*-�����O?��MP���E,j��,��Z��F����}��I���\��"a' JB�4��R�',T��T�ћ<V�@S���ϸ	��iFD�﹩/H�`wz��/�@ِ��ર�\T����#�z�9�5�M��7�"�`��#	�Z?�Ӑo���L��(%�-3��V�@��#qH�'۱&O;���9��v���7>{i������z���jy*���"_l>�nBS(��\w�:�Լ�-�&��}���g����-�-{
�Z���H���@=K�H�������r&�X���������5���W0�@�&	�l���`����U�@�&[����	���۵���V��T��e'_t�}�Gߗ#m{U��Ұ�--G�?��V�鸲�5Y~�y��Q�@���'嗒��:�#:M�"��+��Q��k��uD(�C��<���e�_ϋZr���$� �M�_���F��}+�_z#�w��8B-��aڤC��$�%��V>�XȪUF&���5��&X	����J�C�)�=��ݟB͢ԥ��Z����S��"�FJ�t23?�NnLuB��͆���[��!��h�'\��h�O�$Ꞧ�����3���/���<��?�)��i�mj(S���0_�6�Jw�Y�m+E��@�FL� W�i�Y!�a��d�F�w[�sZ����;{�,��q#ԝ�E��R��.U��K�h�4��L\�>��o�j�--j+���QF�7Eu��H��Jjm}��<=p���f���zZ�����G�IZ���YŸ��¾��C8�&��Y�����OqAl��:��z^��_����t�F3Օ(����� ��5�+R4]�&(�^���̠�/!)�l��
�i��@-����e�����h6�R�չ$�w12^3�1.3}���{kȖ"cU���n����ֶ@XxsX����(J���U�=}��ĝ"���������:�{��H�ܕ6��?���t�2�Y�"���� I	�����D�
!���9F����T+xf?U�tX�mL>�(�#	�++�L��2H��+Q�l����i�����e�7�T{9Z`We�ݽMF:s?}�w}sS=5��}���%ϡ�������� iԂ���V��l��7�(�|�	(������a)���J�L����MK����7�0h�b���Qa:z.Ś����
�!<.m�q\	iJw���8���(1r�a���>姊�	I򼉠T���X�����W1.�7��u�u=��o�-\a�I�\R]�=ˠ�L�� a��v��ЌM�ż�Fm��c��@^ �,S.`�G2��P�>�YI�̢�<�پ�*	vK'�#�r��� �+��/R솉Q*D�I�q�\6�&�Ʊm���}$ٞQzH�K������ENt���挭�3����$-��]2�~�(����Tz�BZ��h�οt��'ԯ�8ϼ\�xz��X��`|��IJ}]�v���s�h������ojf��^]�u�-���p�u^֞L�|�����
RrN|��}�%'&�u%�6:�((�I��n�$�n��K�'-W#��6�d���o4Q���NW'`^��`�M�M�A��00�,/<��xc��7�j|����*��iK�5Z d�� _$���Lȣ:ޘ�������;����x��0�hlġ�]�p`����0/*<)��3�iW��בU�]�W��5�F�:�V���'�x�/tT ��[y89��nѓ��w�X�9����|��*�kH���g�^�W`G�ђ�[x<C�v�d�vU���� ����<�%Ƽ���N�J�R��X��
i��f�����ɏ�&'��뺡�D�?}sh����{Y����2f�{)�E6��l����A$�Ni��.��Q�S8�a��T���&i����0�п-A��̂x��8
�<o[�N���S�.�S���#ɮ����|ƭ[N�$��gz!�\!W�ˮ��1H39?����yq䠅�{Q�ƨ�c��ib�g��V!�A�$�䨋Dg����}߱9�`����}�Q<<=��lÆɦx�U�i� ����;�HK�.��ה�î�_vB_`
�d��L��{�9���M�X�$�u���(k�A)�r��������"�� �ʇ �F�˫l8�!�+~V؞�]gP���+i���i���an2���մ�cu\D���xY�0!��̗@m|���l�݀8D[:wo�qݲ�kKWA��;����{�/i���A��rhʥ�!R�H���/lP��s9��F �gڜ�ӕ<�R|afC��pn��>�.A!�S��kh�i8����U���H}�
�2b�a}e�i	��Llr!>U�)����)��_E���Rڑ��)^(s��8d;k�2JdcK�x}�̲!s2b�E.���P�ݖ��J� \"�@�"�_;���b̻��~Ko/��D�ۈ�zV����.���c���hp�%�	�_J��ӿ�}�6L=��9���i4��	�*�����{��ӵ�P��7�L9v�p���"������mw��kQ
�ص4����^�ݯ��y��z�� �^n�;���<q�c�C�@/(����pX�y������� �^�`ߩ�V��>�
2�-��$i���Q��"��n��z�9��N^�>󥶻i�2�����d��3�ꥹ4������3|�!�b����=�H�K>��"�� ��DN�08�@8Rx�r��9��SϹs��!4�R�x�+���j�姛 �%��f
�<Ho{��߲�z;��CbGw��B�EX�&Pо����� ��N��M�	��I��7��)O�^�d�ufJ�L`���Ao��._�LSZ�$�߈"�]���Y�F�0W�MD�$���bM``Ϗ�B�K�+g��x�� ��p� ���{��W��c�����IXL���xδQ����t�j�f��h�s�9��O >�ƕ1#��M?5��� ��Wk��H|��U ��dswGi��	IwN���%��z�e����8�_���/F�Kؔl���ov�JN�Ҿp(3�-�`��#%�����ۈUV�<�������fr�B��\�`�)��/��� #'�xM�`$���{ `��PQ���gG��kvbJ�2T�I���w�B�f�`���%�!�h��!��$�Z���ǧ���( ��3x�ak��#-lū�#�Z�v��Þ�R��y��L�br��"�j��O���X�7 #���:�V��7[��
�Xm>��*p*�g�t�G*�W7}�SZ��i.MD�O	�n��$�&�2�B�9t�=��&����`����ݿm�`k1���B˾Z�*e%��N�7,���&�r�I�l����F'��C^�)#�yeRҋ-�;ا]�?$��k��Ӥ���2L���ai(2ۍ�Y�ȯ�~[=�ኦE�Y�h
d�/\̹��6T��o�>ꢁ�Q,)3�v�T=�f�]���c�������6��ߋonJ��cVwL���y�_�0Ml�3a�����P�a�Ʋ"��0�yW�=���C��A�E��� T\J?�ߤ{Wm�\#^�:nJ��]���/�h�I���*�7��C@Q��|�����}��3>�q��7�������0ȥ R��t*��I��P��x8��q��)h��ڐ�~Q��!���:j�.����	�G����w�!��W�PV[�`�"�Ʋ�d+���
J�,}�ր8��(Y�~3��?���5�_�Ie0j������!��-~�*2�0\�ŇX©�Ӟ�'I:������ϒ���esUnfM�?Q� &�	���_R?�:ǲ2���fE42�$�Ɉg>�}�f=�_�ҰY�*T=�}�{*b�+�؛]��Y|�?��;�H��6�����NcI��q����	W;�ļ�� DK-�l9r�g"l��k�"�?��V��SЋ���e��ٖDك�J�D,�{X��eD{^��M�9"��&�m�oM'����·M�̿��d4jt��1��O���@��zx�AD���Dep2֋�qׅ�d�6�� ���ZAa]��|�v���l/5w�����*�j�h�oX댝$쥈UQ	�2�ΐQ�>�7�6�72�·������5�ѧ��4��l�"eKm���4(��,�����p% >�����p`m��U��vZO����6�ft<��ܒ�$D&�܈úќ�q��=����{��r��~��_�E���`x�FH +=�\2,]V�\�� ��V�a`���=��yyeIdr�j_��g>�Rl^mpZG��`�D�3~п�b�2����8ڵxJR�����N��z�5�?^�S�V#\�1y�z��YOI����N�#t�ӄh�Ѧ�tpt��{$R�d7�.����:��u���ǁps�/1����0tm��+s{"��4Fe�t�O��tL�Yy�i�: ��kj�����YW`l�k$�;�U��	5����f��,�<p7�����X�� ��V�B@�U��A+�3d@0J闎�{���;�����	��\�,��Z�TG�%���"$�������q�������	U7�8-R��GU}?6�]/���&��?X<=�3���1�����G��ΑSy��[�AXܨ��V�����m_���q]���{t#����r8ؖ��	mү�70���FZ����Gn��>I��64����S�_ޗ�����yg�b��jV�/lՃ���1 �"����S��WPgI$A:�U~�Ŏ�~���ح�ٿ��ՙ�AQ����Q#[���/�'��l\�w@䬾��1c�i� ����r0/E,ˡ�>��͇�͞|��~��f��D'5F����u�7jEO����z ��Y����}n����I��I�USxQ#��:q��x.�啂��8���
�8�G�`�_Ʋ�k-�����I�+�".Q� 	�=�@����%~���kLG��`��E��nI���lw��%�R۳8�Γ��%Hnِ���9*Y�D'd�	BQ��z�B��5��K��N��k�%z(��b�88������)�r^�<Pw~g�l����"�-�lf�)(��f�*�J8��4�);"�[��֏� I5��J �ŝD�TȮR�m#�,�OS��M��cJ�mh�wY%tW�~Cx���	�B���A�h	�g;� }7J7�TWt�t�Ʊڀ�O����/�ʂ�E��_%�f�(�u��+������&�R���/�q��A������ZU�؇%m�H�'[���Jw�e9!���`V;�39����V*" �r#���9�{��I�@5���¼܏,u�©*D%�!�G�e����0�vX�R�_�ʦ┍hG�r���W����J����F?����3 �xW�l:�I��#�d��K���1�_��t���V*J
�B;���Dt�L>�UjWso�V|JA��x	��M}8r����r�?T�_����P��!���$O�lr~`�#g���L�*.g��2Y𷶷fje���%��b|fzwX�Q���ҝ���X�A�Pc�'�xOt�?�Q�л�E�ٶ�?��DY;�tn�Qe�����`2�y<�t�����G����M�r��#�<R�$�h�|����P�c��M�"<��d�'EC��^�L���:3����Q��^���q+y�Aɣ���?=7둯|\�03��(I��P�`�l�^QL���`�Rj�N���2�Z�0��S(���Bɞ]����W�l�;!V��c:�����A^���d10�9<G�T�M^�1Y���L�[��ȠT�>_�X��s:�j��W}I�p8.��P�}�쯇�Ƶ�R�XWh��������D���tw��-�կ�H�A.S�'��U09�Y���4(;6���ρU��ø�g��U����ß��'��I�k�Bӹ�-�uo:�l�9���ω�"ZJ|-3FlE�BH>���ȢPX�E��<�����pM`Ŏ֠�z�p4H#"�Eֶc>X�Ĝ�����So�'���9`X�d��S1K�!�a*Ěl�M�]�	�����iaH6-�?����O[_��i.���@v�"ీ�/܉��xd8��Hy�crC�j4�K�U�B��T����"��*?$���z�Z��u���	��.߬��팊��4�%)�wE4~���{�&��m��$��ڊ��N��oў t��O�_	T%94�8-H_���J_5h��9�Rp*�v&R:�,�/��
�[�^H=1(9�w��/ ��H$at��C�����9Zp�I�{�SG7�h"� 7�.q[=��D�1b�-�p�;�(�����QT��Ϲa'�9�TTy��! M̟����;���`����s͍p�v`~����>N��N�f��0�Y�f��r3�ָ~)w�QBAȃs*z��޿�{ΥG\3=����"&�FJ��ϦP��ˊy������p�_U'q��j�%��|����m��������E>I�cp��}#�h��B���������=�@�O/�bԅ�Q7ڵr��P�Κ��>���:~;<�B'�
r���rr��bm������
��1�z�S�SoɿV[� `��K�O�7G*�8����.
�o�G��I�9��r(�S����}�<��)m��]��L�]\�~Q�u�wc�k6�T��]jk�xӴ2z������@@!��8��EԘW�-��4F��)�n��� ��W�Nf*{�*�*U��V�^']$ۦ�PE}�q��Ub�w�꒪���/�{�S�嫢�~���B����Q�@۱��t�'d՗��*��5:4u�����H��)h<@�43�*��5:r��?S��O1������I��x0��� Rn���C��g��7ztWĄ�\P��e|Gmw&'5��Qe)_�5!}�t �$.c܏�c^�ibZU���T拶��O��5H��V.��t����GR�����0����:J�L��0Zk�"��w�\b)���;��/$~�c9�X�˚VC��R7_�q�DO_�itΦȆy#i��� ��� �J�T���ӫTJmPn�7&��֊�s�`��G�ؼ����Y��E��?�k�d�/-�߄F6�<�g\�h��~�q?aAs�cjm��j涴�`�U}�М�����ײ�Wi�O���TǊHu����0~18�Wܧ*�wZ�u��d�_h�-
S����W��p�h']�Ge<ٜ#ĽQ�k>�A��2��.�Љ`�|\�"A`��Y��mA?o|��V���C�q��?���NX���K�$yIq�g�
#���	l�O��n��0����Z�C�`�_ݠ����K�ӆ��������g\`-u���F��ڶ��nZ�p�4�	*e��w�u�m���@e��Lw���@,�x"�HX�t�o(M�gͤ?�]�/u�{i�=�����U
]j6�M���jrW��^�3۶lי��{ ��0s���D�F$����R	+������@'�MĊ�I��"T��2�3�,i�D�P�ldj�l ���L��V����՘�  �,s���LGӼ����p���|�A���A���WY�z�"@ɗ�~L'� �B�-�r���Tމ0#ڶWo��GS�>u/{/
	�y��6v��۫C/�)o*��&��t�g�(�~����Z����>r�Br�}{V	9�s/���^��u�C��BOytF'��ϊ�<�?���bT�%�W���pӇ,�dr4���0����>�w���	=/���S�Nu\�x�e��v�̒��Mz3��?#�U��4�>J��V9�N�-[����.����TK%���B���+�+�4$������� �H���Kbl"�|&��}��)l"��h���Il�Z�H���-�Z�.����"��t��0~�l�˃�7�ũ��9�fڴ���Z�5&��ۻLW��?��z\�K�74C��z�̺�j'w7	ԈG�ŗ1+��=��`�x�(�'�ʸk�@V�i6�]��y�ٓ����hodPn��k����7 "K�������}���Xl�X�ۘK���/*��Y5vzA~�M	�Y��u{��Յ�ۨ���izm�y��B�9+AX;K�ݪ�d0�E���h �������b��J��|�� �x�?y#wo�{
�Z딐9��y��Ϸ�4�� t�>�&��@�'�,x�:j�����i2�ī����Fp�9�Q�%��""������.ͦ��7>�n�p�܌�yk�}�ޛ}�ۈڤnB��Mx�9I �Ėe@�����A��O0eo��8e�]��]q	r�վ�U��?��>�7��7�7�&ȼ4`!���&M���V@�$;>lt�~�������a�Z��eD��M�M7=�0
�M�j�%����J�K��A����d�s#�$ج���Dm�5���	P$P�Ia�����}�����������P��z/u���TH,�m� 1�NqK��vr�,p��m�ǆ.���j����Ũ�M[��K�[G�[�⊁�==�3U߱�w��f�lq)��  ¨���+�wq��+qf{&CAz�]F�հ�%��~� �}5P��I�{�:\������I��\����$N�p��|	�/�y�Y��4g��Φ�z�{�m�Qa��F[QUO"?hk#G��ց����O�a�s��Ԟ�
Z"x�\��rЗt�
J�7��L)���T��R/e���*�Beo��;��6d�(r�%�Dy�0~B})�h�g]�˶#]:���4Ļ��16���b,|� yȁ�F^f�]#�k��fH�������䦗�����H�����шcԑ���/c�C���z-��^H�$��y@���\{���n�^��$8�~|����MW�:S�_|��m��J�vP!���0�J��`j�E�9JV������4��\!uZW*bt�O2���e}��Ö'"q�W@3����a0� ͉���fS�]��s'7�jA���Vp�b;��h�����g�i�.ח���n�Og[����K_S���7M�K�H,1�~V����i7�C.$C���p�,��ZZ���� �Rpn<�=��9Y+f's�l�DO��;��Kx2\`R�z��z�2��z=�Vd�G^Q�tS{�oL�	�R���#��dN^60����H���A��-$�%'��(��EY)t*�� }�ē�F���:�GЪݪV���_Qa��T����l�M^#��Z�B�����{�M����@1$�'C15W5w�ؘ���La/1>�W�o5a;��t5I5zܖ���)_%���zj�%��6G�t��!�ц��]k�bC N���#Ѩ�7[`q��ɭe"�DǝT�;���`ka=M"�$�
ԲE�3�q��0̆�G4�E�c�ڣy֖�F���3I��N�Kk�&���H��:1B�;8�:���,�*���â����̟+�B<��F2P���~�P�N�W(A1;*H>�X����W�|rۉ���,q�����������&���C(��,���5�T�2ӛ.��֡�
e�>Ӭ�V���4�e�ǀu�s���PR��+�԰#��J�Q|(�
�2
���L��?Ub�*՗�ܘ����eα�+�U��Z6����I=`�d��ٿ���j즜S%�W�c���э�@}Q�y����@�a���v�{�A*y 5�D���t"�06�#<Lb��I�q� ��h�l�` �o�AlAp�S�l�t�"��j|yb�ț 	s��=l
v3�8㱪�,HS�\�Ir�KCa��pz"���s�9�����J(��������1F�N��N��J����~�����teq4�|���`�<�(�`L�\
S�	����o)xn.���
1�͈��ѾD��7�լ�+l�m�L��Cf��O8����y��I&� 㫖ZΫ�\�4:F~���B� ���Gy�^��f�4D�qF��$F5�G��t�)EHN�Vbw/���Ǧ $zh����嗄lbGWp����=%�����Z��i�\t�7��#	�nۀ�aB��m8F���D�ƹ�qerdr=���~�Z�quϝS�s�x^��A��M�G�g]���� �ΔT*�H�0tvN,{]GQ�#Nº��i�vRQ��׹<RE�bN���f�z.|p�?8�U����WW�	P�����>ъ������^('kym���G��kB�K���
0�A(�,��=��n�w$h��4���{�_"�-�Lh?����m2v��U�� �u�"n0Ŗ���U�p�V>��w$_q8��@��T �)���@3��3��n�-��7��*$�n�V���=�{!���Gs������g/�Z9���� �Ϸ���܁���3e�y�]gC���w���72ܥ�FdIp '�I��9!�쓥�m��F\t����Wvn�	���0!�I��Y}�*ٱ����$Z,�w�7��т��5�~��V��!|�d(��,�N c�laX��s2I�ia9[}����=�Ф�hA��^z��/P��Z�]�m�3�~m������`�҅�j��r_�[���WEr�f�.�8,�ܫ�Hw�|��!�`!��Fg���H�%���ǁ�2��@�Xɨhc'�SJ�5�l��Ȭ���_d�G��\=�(�V���3�j-����e�P��v��~���x8]�Q���[�P�Wx���e»�������֩D�����r���.gu�Ń��(��i@�i�³��#�E����_^#%M`�u�4ru,f��	���ϤR�)N�x{r6E ��ӯĽP����.cE#Q���d����L�_�k���ct��|��3M�����}������9��@�k`���h��p�yf����K�7���4`����:vVOR��vSJĉ���Ȗ�e/$yhy�F��%�<T�1h�f�����[#2лӊ�(~3[.T��?�N�%N�%�)�N�L�ʧdU>����}�%U0��˛��;P�(Q֫�7�z���*}r�~pe���Le��'荽�vf� �F�k��Ƽ�ڠP����"V���C/�F���ل���O.E���,G�N�e�D�f�������gR���Ɛ��P�~R���l�&-��5ւ��d�Y��c��tp���]=D�=�����YB;Eab�~]��^'
�^'t_���,���(�0�eyPD�~0�fQ�s��
#R�=fJ��I|fɂ;��0i������1M�1Ϣ2���&��8����p[Ȝ�y�o�s#��s-�St��]��e��q�(�`N�"��4�9!�~��Q�-Q"u ��%��^�!#o���O���Uѷ��-g��ߥl2�YrEnE<~-[:�p�>�Y��2(R���{$���D�|K�\�Ϯ�֚��X�7+���C�J�������1�?{��No��+��S� �;�BLVe�1*�e��]uM��Q�G�o�{7�M�5��o7���N��H�������J�F���ZQ��� ��t���~������o�#�G����dYF��ئ-��=pw`N�K�����C��6Crc�O9z����k~*+�� �[�������znR��a�1�6M0�g�1~k��t)+ȅF5��#�G�m�./�\���iL_��$H����E5���k� o������Nh6T~iV 	��Ћq�q��p��W�/y������3�Z��6?Ŭ�>��S��=^ΤE���� ��AL-t�4�O���v{j?`a��Q�ǖ���i.Q	dfX�����ߡJB.�w��_�y%7phD
�p3��F�A�|±�u���Ek�R1���T�qkGɤ�\9o۪\ӱcN�=rg�nt{���@�Q��KRG40�c`�Zg�V�nd�x.��J2N7'r�'�L�5�p�F��b��'��^-z����(�%t���d��̱v�F&Q��+F$���szL�W�D��
����t���E��H(a�h���Ӊ� aW�%��*�If��,^��I�c��ޙ��cpe�{4}e���Wm����(-�(|X!�l��p��_���t��̾P���j�=�W���
��8�+��V�2v�~�sd�����N�Oe�<x�:l�`c~ժ��.�^>�py!G�K�	�aI {����6!���6�7�!**�C>+;^�DR>&U�Ta�ni�p|׶�����@!9�����l���y��|�:[(��	I���, (q�#E�A^���2�Ȣb�waw��{!ģ�1x5n��A����5�#�}|B?���x�%�+�x��Abs+�aCNT``�$��'���V�gS�n�a{u����o�G��j�Tmb
�-�k��IMA���d�}wS:�z���`�&�{h�a�>E��Oٷ<�'���۩(,�!�~����$�(�He����'e�\��/�,R����S�n��Ë��-u�89�[S��:�
����/�U/L����a��S�H�M|?�C�c�0^5"���0g�SK���&.oy����B#l�qT�x)6��Vn6���;Bz�S��_L�`�l+]%E���fAe�^�DыQq+�g�}�?�jl�	�H���0����k����r5#�d�v��<BF 2,.���]Cf�������1�aN|�a"Xc��qī}��.��g����0J�t�t��*��,Nr���Gi�_-������v�ׇ�VX����U0����%��42���]J�;5Q
pC��M����1�`R�T�T��t$�k4����Q*K>�	�sc��޽%=vomO��g�	�i/�^�b�x�:�A}�^̖9~Xc������q^��%���A}|���FF���?ÂOR�4��F�R�3k{�&�&n�t�H�ϸ~����}�B�V (]�$���\�S�j5Y?�`>��$�s;[|����U,��n��J�Z�$�dh(�WXa�Y_w��a����a�L'Uo8	�(}L]#>|c]P��>Y�����+���*oG��E�!��w'�G��T���`g"�ט�1sj!hk2o�jEF�2�m���g2�B�U1"���H�2qd�� �&P'�9�u��5%,�25�^�g0�M�_��\�I�gn����0¬�����^�~t�,�g�$��^*y���x���xR���}~m�0��Y�?.��ӆ��e4skI-~��	�������иO�4�?5M�QZ���uPp�bKK��Bl�ʼ+	��:?���Ǔf�s@Hu���E�Ume߳�B��=���P{����ən��hΕF�Elq�~8���߇�؛X|�t_B�<�o�_�ޥ4�Ղ��lkMУ��O�,}R׸�A ����P��X��}y��o9�9 ����u���[K"�ED�/[�7�� 8A�,Q���-���{���	�Bc{��J��������ǀ�(/��
�T`9:xw��i�R�Ù� V�B
��G��m�l��фgs�2��*��
#�z\��&��*��}82�pə�E��L����=����� Wvq��秣�FTs���B*�9n�0�,�̤3�-a��YL:��Wҏ@�����NgO�IBPץYdG3B���B��)3�B����Ϋ�fAM��*J���A'T=5�bo%�B�q�%��� !�C�rώ_jL�Ӹj+L:���-[Ix�$�����Hkmt�Y��C9\��.���2� 
��ʗC��\�M�kΖ�wo�)��u����c���f����8�2���K��Oh�JGh�����_��	����G��������w,9� ��&O]c�r������-�ger��a���i���+"Imjge6��q�Y�9�|�g+慬;�q5	r�R�;aїQ&}�����S�L�:��=��I�S{���I��4���*0V�vpJ��$/nL�w��nī ��O=���R��տLOm��>>���2��%��7�U���u1�����_�������L�+�3}�Ҵ;�������N���'!(HX6�Ea��m��t�G�0�������џj"���ǖ�7��K�>F@�e�Z�z�Z���4n+�Ř4�l��4�̎��1,H�Pd"�;<���r Z�~��_Ab\�(�m�*:x��a��囦!�� �4ܯ޵�y	~�*H.� �r��q�]��pI�Ժ��ǋ�0�[n�a�q��g�싆Q��9�r"�_4"��|(��s�H�a�0E6�v�@{�Z���TYx.c4���)���S���;�1��y�-�S�� I���Y�y���!�UM��G��#偒�s>V�Q ��ԎTx�v�O7�t�	�e�z�`��6���n�R���h��G�=Gp.�^�8��?��cs���6��nN�t�6���~pj�a=�"�>�Yy����p�MZm'i�V�)�.��]�'�1Ҫ���t�SԵoRK��b�#�~]=�'�����|�,��䵈z���jDb�\Z���f����+(��v#��O��כ����߀�L�;ͫl3���*B �����r�A���22_Գ
�nm�����l��(87(70ښ��I���Pۥ�	<�[z_yJ^YJ����z�9dw�� �$����L�U&K�-;Y��>S�Q��߆ٞ����?p{0$�ԭ��Mfbki��i�ĥb�a�.��?�[��ҲC�Љ��%�+��ث�\x�AI���"}H.i��*$t����5��ܑHa=�6L*���ڪ���3��88��E�?��A���.��U��^8:�oprk)��rI���
=L���Y����ׅ�P��T�^$�� �Y��!iő[���9�w���Q��A��E��}=��:���9_uGDJ��#0�������`n7�S��`�*�w�b�	oR�z�ҳiڄ"��P]��_�"�4k,l#䅦�lZ��l�	U����	\�Q6����7x����!�-�,U�_(q9J����=[�3YFF�r��O�yi�]Q�:�z2BQ`C�[���6�H(��4fq��E�7m���s���h��Uo�n��8-�ꥣ,��g�J�bxO�C�P���³��v	��Oty���&�]���P�&�#��x��&kA6���N/�a��w&��PFHTra�L��N�c#>���0m��]�Q�z��v��b�T�F��7�9i��a��t�j��>P��n	�SC3�B���6�L��ә�nG�U���]�RiQqu/`]�brG�n�ܹ����v}�E;%Bǳ��殄ms$x�8�vgU+#�ђ4~���e�Cg��](���f�z,+���U�#�Ŀ�	��N������ǡ���VOJ!�>�NoEV%�`�>���iY�݃f�zE��R -��hI�͒�3)���T��״p
��D���p\�mk����f��cʸ�l�z#Qu.�@�)SDE�o�	�4�y��'Հ���d���8%mO�X3e�T�%o��g�c��f 	�%��ƛ��0���B���C��;O�fM�X�����{�T�����?��8]#i|����Ds����1���O��C��ϥDٔ),�#)������3_v�����q����(S�r��0q5���x9��}��c��2x��\K����} �@X�=IHUF���4�ݺ<��x7�-i9���:�ٸ�,<�Q�`�Uk^�;m�� �������E�?�뺴����n��X�b,K1M�������J,�wʒ>�C�笾xEژ�_���,�!�h�AxڬjԦm� ���K��2ES�)i��N�J�a�����8��p\Yֆ;�v��\�i��X?M���qJHq� �����}O�7���Il{��@�3�ڹ"Z�A=��"���6���]A6�dE��m���璉��,b���ڠӍ�!@Ka���G���9V��C�}�:��� ,�ϭ��[0 sz� ��oJϪ��-j���>�d�����(ť�a8������7b����y�+�/
�ߔx�#�3�)@�2Ѯ6'U4��dס���7�S�ldפ�ȩ1�w��78� ��b^����:��~i�e{��B���ľ;&i���9M�QmQ�9���z����C�J϶�o�u��"R�TO)���Xp��ϣ����"?�eW���Fm&p9�?q��g�r:*���sm�$G�\��@�S��0��/rh��Y���D�3�s�Q�!�Z���F%e����LDvջ^��f�h�,88�����G�ƽl�;��qY�-���Cp3}�n�?�#���O)�����V���W	��0)�L'�68z��L#J�p^�`��w\��KI[���t�n�<
"�9�p��#d�c�f�����}�	W��9JT������q�ݛ�W�T��<l��T�o����ЎE�ӗ���S�V�W��a��X�s�2��?�����=�x�J�1x����k�?B	[����? �3�U������u�#E�1�·��D�<�c@�>����dS��F�~6f6
$A�ķ������N�r��YQ`��]�I��<n]@҅��<�c!��6� �Ly ��N̑�Wg�}��&��W�,
� W���i��D�1CY�F�nGa犇m�լ���}	A��p̆���ɼ�����i'��C �鷱?�%���P'{�df5�j�s��q�ns@��9+m�u{�7�N;��6��\%iEh@�ͫf����)����SWܫj�!�Q��vk�x z�D�; P��,nVvxXG��W����@��xx{{��c=a�	g8���t7���W����rp�u�yl?N�<�gd�Ygn�5��^g%8e��lez��1�����[t��u?���5��G����Ґy!x'�zn��r͆	����_"v�C�6�s����LOH~@w��;��l�@G��*j����]__+
���{�QL�ċ :��O�������Y~р��rT�ĝhȻ�����L_��7�N���D����@�2��r�aG=�xO�L�5��)�$��5�激�Qm��o�JUY�/V�?�����	%	�gv�QB��r��zK��Ǹ�p:h�>m&�;�'��qF�3=a�ߥ�;%Nvx����9�]��G:��ޛk�a�Bp��g:�~pX�M��Ww�&�,�"'X{�)���6^:{v����4%W�Bb���&�� ��H�}����g{H� ����Uۙ���?� ��Ӗ���83K'�k�G��*��y���q[C0��+,YHc�_ V�&���7����W�A���y㢝�nuQYl�{t[{��|K8��}]*�1KX�y%ަq�:4*~�͟Fx���EU�P�o�tS�&���&ԭ�zЯ���HV�/��4�=�s����tM���z[Y/#�3�g�%��𥙀BbnAL}����AY:���w>P����s��ٍ�1/���P�A?9���A�Z��M�%Z�C5�2o���1b�!w-YT����9�3�p�1�)��� �TH�����'tH�"�0�!�!M��}K��>��2����8����Y��y�&�@sx���r��@϶��)�~�9Fw��R#�LGT�dJ���,H�l��9z��lY��.˓�$eD��f��Y'��N"���tBF�B�@շ�1IS�HxSd�j��=�2����|�$J����M<������m#��Z%b�_H�B��#@@>�6�um�8GW�s/��+�,�ҏk-G��o���&�ig̽�<7��0
����݄�?�Ԥ�b30�Y� �mx�j���
�#�/c�����7����̛3qa��L׻r<j��5�US��@y@����\��j�4s"_#�J��A�?W7�!�w4L$4�	��tO�?iC�_�D����d����٬����F�y˰�� ����i$#d��9#��p�`[�Ky�,���MYjVg�/�Ic��������8���9�b�RR0?�mb�8R��~�旘n�̵)t�?�~^��?KF2oH<,cSgK�W,ޥ2�AN�n�f���e�M�%��,�c+ʑ�.� ���(�ͬ54���Ɛj"-av$%ז�eO���q��(t�K�
�*δ�A��9����
�T9J�~<}F:(�[�F%���dP��v�]#�sw��V�����R��9w	���ﬆ�Fd1AO����p��Fb���������Y�����њ���
9�ؙ������D�\����z�@��*� q[�[g�e�l��#��`j?@�-l]O�;��,����-{��œ���s�9��;`�5��ްP���O��'� ۦ?l��r�����u�����I�_u�����Hߵ���ɡ/�N��p��H�՟��yo� e=�a*�"!�%l�Ku��}�DA�*B3���C�hO}r�/���#>�"��Q��	1�Sb�:���L�9C�';e����~�&��%>e�{���gaĺZ�f<T�(_���Sn��&��[�i�'��'�k�'�Hi��{��6qXSg@�p�߸<�Y��1�q�]_,|O�q=)�ٶgS>�ob��z�
I��u'
`����`�;
�����D�]�{��jo��wȁ�(��{�d�Y��#�A��A�ɢ~�'�P)��IE)��ź�59�,�>V�HA��M�)bh��ueU��>�)��a�[�
_�ǔϴ� ����ʎ�n��FlIK��V�d���ۻ���VQ�����H�]�v\e��� 5D.P��j�ˤ��7ɡe���y����&��\ZP��iY��ƽW�A���4�(�-��+ŋ�0�x���������wY�}�
�\�+q�Hc`(����Za%�_�ڑ!�N�d���b��	��R���8�$�+��w	���<C���~k�i�3~% �S����9ڤ����I43Z@�y������g�v��,V.]?��I�g�w�x+7��;�Z���@��-�j���Y-�c�$jy8� �fN�ym�\1}�N8��ũ/�t�#��+G�}[x!p�ŌR��������g(���ȓ�Ȕo��K�f%i5\i����ۙa�Ԝ=�tk�:w�A�Hq�]8_X�k/3󥴚�L�o�K����#��	;�����􇖑�	����ٙ9"Sк�>LL��z�r���f�G	���H|���U�?��_Yy���E�@a'��_J�C����^���%�qٞȌ���ͤ�q�3!�π�ٙ�t S���uy�5NM>:]1��.xw҆���4�@�I��v%�8�%w!)���Ǥ[B��e���L�\��\/5y�����I�@b�z̔��c��7�Rs1���Jr?k��,��R��[@F8$9���ʬ�jε��LDq��=��?�$2�ǉ�W�uN�6�d����^�|����*Ԋ�0r�q`�z���,7��X	g04R*�\�D�ISm4��
h��Ņ,w�4:���XP�\��B3C}��p7SN��v�c�B�P# �$J]��s���@@��R�õ)�^�� �f-(B�՞?�S��D^���t��<�S�޵  ZR�$2��Z��ߑ��i�Ǯ��P*/�FJ�ɺ���0��$�<+��F�ʩ�s��쓌��w�qE@��Ly�{��rKѓ	f��k���Y�JʎGZ��xf����5��&E�`&ވ�G�锘bˀ�����L��Yg��G����Ӫ̏i��>$��XL�T/5��Ɔ�؆V��m5q����wA�W����D�^r�{�"��(?�f���h�͋�nj����㤞���*��].�dq����x\�÷"5�R�]�E��K	^��xb9���^�ڷ#a��S�#��U=����0~�F�.֯�2�n�i���W�����j��<�#�!v猨���7tݞ��X�!{ca�a�$NI褏<4�_-<�������~�״J��c`��!>ty�h0�-�&\��d�e@����gS�W�?j�=���au��O�&���X�qi���a�?�ӄPU��b�/��hh�hxY|\{��Rk����CZU>�7����<H�0�*͜��²j{����S�u67^iLu3�ގ����h�柳���ᓽq��0{g�$�|�h,�G����`1�Z�(.-ƥ��$^�y�����ۧ
����"���b]�A��P��
�!��NԷ�_�s�m�a�	�@�����D�_�D��]!+�Z��r�1h'�g�K�łf��n�l'b3zT�D$��0w�}�]��,#�I�]��*	�	��i�P���ݻ6�d-�Z��x�͋�W��c&��`����ȵ����Y����µ���GC��k� 1'TA�7������g��Y��(�\����vdC�Y�����)-� �(H�
 ��1�����7б�<�9�N ��BU�{:���0�����Po�rtVĀT���h��}�2�YYRw����3<\���n�רT[�l��R*����+J��=��Q���ʆˡ�S$��я��U,UH�gܛ�X��R6����O��;G�*�=E�ɦ���P��{�%cj�y��gǤ��� n�]�!����z�[���Y�oSBe�@(v�@��:����+�NѨs�K�*{��@��A8����X+�C0e�,x��WY�&��x(X#���~���-`f�]0�w%���Z��L��S�IF��[}MD[+�g`oahJ�R��q�k����iM"�/t؍?8���c8�@&d�P��,�?B�"L;�9� sv�R�$�I�>w.���}ްT�q��ׇF�Z��Y�
�5;�Mz��L�t����Fe.u�������Q��M����e|�s��j�OE��Qb��=�?������7�;���C��,��U\���ƿ/�-,ap.!ʌ�E�� ��D��+�M6{YM��]:'{
M���{/�q=)�w�� ,">^#I��'���y�c�i	�gґ�j�l+�s�d��`^	�<L�H5����e�����*�Eta��g��5Kq�1[��2vw�	��gT*/9��m�.�S��UX�� �+`� �A�Fk)�4_lB��xgl_]A�Cޣj� Za�(Y�_'��MR=���msj Gc���>h`�ێSjc��Z1���~l�O�!��0����G��Ϋ0"��� p�K��ћ���/�[�'�C�A�������v׶�d�o�.'jc���(�i��!�:�v
��p]E��3���4�� 6��H��(�ֵ�B�C`Uz5EbU�B?!��ָ��>��<��!����l��e�WO��f ����f�j�
�g�[X.�4�&7�n��}��E���,'5��6��&�:��T�`�,��|�3�X*ө}��m�AUy0����(��v�N��dnN!۳R�2�
5T��^�����g����p���KXJ)�ٔ�9/50��!��5mIN�3�1���Xj �P�s�'�f���Í�����A"�2@�4}��7�6B�K'M������3Q�X�x�Y-�h�z�j�5�����
�΋���m�ޠm�o�r�k!������q�N�lӷW�$�\��'~i|	����NÇ���� W$+��K*����j�t/��T��> �V���A�ߕ=���,��"Gd��9�d�`��
��"�]��Bp��s�%4i�j��#X��cV�[/B�6���^��������O����;�8���ڳ���UXr^z�^i~��	F)��hU���:[_~��Wx�
C|T-B$�`��g���%J�oXe���sn:�U�?����Gd�2�r��:jղ)/;�D�D���s�yM,���L#�{��%(F����>aZP����f�6��?7`�9a�4GF=�@�fR{��jq8���1Q鿰?G1��.L��Ce�n��������}l��x��a�5{�`V��JӚ:�D_���)ک��b͌����W4�W/V��@՝�cY"�`P��ѳ0�����1{?H,-�"h5Bu<bI���#���Ό�u�&��1�9a<��j ^N��ǒ�}��rai���P�̳�F+.i�Pp*�\e��ąC�U������6G��VYf=�ıpVn9��S\�,�SޒF�������y�h�t���R��	6P|'q6���'�N���������]�b�6ȗ�i�>��ͮ$op�=vp:�5�$����A�ƍb��J[j���¹�B�a� �n�4�O�Gx�� O��+em�n$�w�!�/õCh��i���M|�$��� t�/��'�=���_�4Rm3�Q��<�aٍz+�{��6�|�6	۝{dEd�w�A�b@������ �/5�p�,5=Ԍ��T�pR�F�KMe��j�����n��s���&���P�����ȡ���W�Z�IIE��	�.:i�@*E2�����u����:���S9<%s{����_�k�W�{�[Ȕ!�PJ��zT�vXh�X�D[�=/&/�!L�&��O��Q��?O����&����@���	'�T��m�^���v�$�Nׂp@�0��]�_�G��]L�<%���"]�Lz�j�����H(�M�^AUC���3�g����%L�C��kq)���5�lڗ7aj���2���wIE,��c��GF{�tg��	�P�7��F*�"�Ϊ�Sٿ��чD� ��GSSԖz�,|W�1�
p'_�k�ﾨ}�6�]a@*��z�Dg��
@��=��V̅)���D�0�C0{:xa�Qt�w��I��E��R$��,�,�ET ����= �S{����~N7d��;p��-i<!MW�0�����M�9�/+O~N�T�E�?i��a��,N�PLgoQw���{�_�v��`����mV� �1���ǔ��P���!��DQ��%���X�k��\�^lb��Mr�M�W�KH-���9��΀��"�vZ��zn�	xQB���V)�Gc咆]��dT�7���ל�e��oTwMױS��2��>����yL[u�\v�ۛ����L*�k�s�o�:��zr҇�5ad
��� $t�J�ԋ�\����"�����=��v��h��u�p��HjX�4�K��e�""'��tSp���0�
f>ICL6����q����0�?.�R����d�]�gΠ��#�]#>�c��]�1�\5#��x�����Q��W�6�zX��� ʧ�x�Ҟ�^�"4,���_�4�U*�{�'R�Sr�^��X`b��6��2Г%Vm��dT7��P�ѐ[�
��*vʶ�Mkz���f�=MC�J_�-?����{P��U���s�MW��k�xUD��^6���6�Y�e���HNx�ɱ�!M�@���,���&�I��b*W�J��������/�c4�����6���v�
Od�u���B�/��*L�-Ѯ���
�;[�K��Y΃L�"Q�74��1, �D�U���Ф[\?�˥?��[,��?��kXi&k���Y��s�жT�E���y�x�s��k`� g\Z�������[�Ut(� �5��L�㩗>�lH����޼���m^�G?~%w���j�	ũH�qV&ӫ-����Ƅ�k�8��h�KVf>#����:�1��gk�W��v��
�ؑ�1�m(M���K�.���EkR'��a7%�`�ȝ�?��u+ �V�:�2�t�H�$;��(�;�T?�k��a��W庸�O��q
e���Ռ��0�� D�L�g ^ƯJNˤ�*��H;[�`	oK�#��M�ѨZ������s�]��㳥�.��f���Q��v�M6e���O�'x�M���(�X�و���@����	�r��h�eC��H�l�[*��i�86з�Qp���{O�n{mL6���U���/��@ �M\�lJ-=N�����ZUj;��ஞ��p�P�G �>�KJ�O�<f̓���̓9�WJ��tun1?����W�3����
j>!R���q $����b�(�@q$Y�ÊϠ�Dߛ����|�F���Д� MQmX u3�K��'HAgj�	��þ/N�R �p��w�>���8-k��]k��h99�f4��'�H7�@���\�~�w(%-kЏ+� ���j�
��YX59\���n���}�#j�|�:�D� @�h�\� ����}�P�o+��Lh���A1�:��J������#~�2�0�+���
/%����Ңi#"*&(�w��F'����zbi(��`Q�����a�X�4�W����\U%0�SO4�ؔ1g�����eF@�b�C�v�Ã��$�艜��8�挰P�? -��cz��R�V���i�i�^2_ˉ��8ro���m�!�:����hNA�aƨ~@�"��ڌG�:�-!��R���u1H�!�*�/>�L�Q��2~���!�����A�*�A4P�6���=�{n�+5:b-���:ݝ<��I1�p��y�!�I<���ߋ����#=�ai#5^�t����)B�DY����i�Ym�����T�`���<aD
�
���ۦv�ެ*go<�y'��6	Qϕ�O=��M�: d%W(���b��-t�\G�k�����P��	��`�/I�<r&�v�K�?��Z����e��SƷQ��W�yU��HZ>���r�5�o�Й8��꫕l�|.#��FT��z�$Kߏ�,)/�? ��aך������>Z
<Pڌ_�U� K�x`���R�gX��n���[`��d�7�W��y�WL5�4e��A��t�ʃ�tM�Q��F,x�#A�Yh�m���淰�5M8�Ӏ���Ą��ǐ���zW��A��K����ڊa�d������I�jY>�q`��gX�3��'N?iC:�GI�0���r��zi��L��@��l��0������}�C��H�������$��rg�)�ˈW�ӛ�^RxW,1��d����zw+dG��BL���	���eO�����U��4��z'�*����³����Ϥ^��%��Ϲ���$�`W�r���j[b�W�C;�3��k�GW�[����e2\��a����԰���;���i�.ȩ�X�F��
C�g)&�#�$ڮ��^�_�ꂚ@�7�D�ڔ��OkճscX���*��6�k��AD⯥���
\�{�Oҁ��A���1Ϙ�V	j�a@(g���$+^�Ml8�}��e>�PV`9�@� T�o�$��
��4�85ɡ�4�,���^�T�]T�+���D���
��b�B@3���2:�[p#,5}$C���!�y�x{T`�H0
1@j��Q6F�\}Ֆ'O�f���:���Z��"�I���	� �����r.݂����M�ی	�u���f��r����`F��S��.jɱ8uR��M�z�>�����#��'�6oB���J��z�ku��;'7�8.�Qs;�T�#E��3;.� ����g_)�ߒ"
��9,g��Ȭf�sOF:��.�S��j�k��n�3��>I;N��3}\��}@l:;��]���C���o�:�x�0Qv��s�K@gJ��K��(P�n�rЏp�o�Xp*�XrX��U�o�hø���&p��m�n�[ALȑ�O�h�2+��dL7�!4O����B�9��h��k�s��_��2���`��)��d�/�j�)�2�EҬcXT"Gw`ILy+D6*�W[G��bM�<6���4Au�c��kO�M��R��4�n<�1�;]�.+֩�aY1?�i�q��kv���q���^�C<�jNB�u�5�mAs�G���.Ј���.�����
�7`���R?�{Hwg�e��酹�c�@8��)�����i[�`>�Q�N�1a���6����X�L6�(�p+��U��-��r��f��14��1z�~���Q�t�%"�r0�ʾ;���S�o�s��Y��]��em�v�wg��\T!|y���o[Z�X[M񻮀�t�m��5�ƏI���ۇA�I��u�J���­���/��u~�eɳ���\�-�px���2��+G(�Ί�j<���;�v�F=�A�]/!ߡ��(�K�R���e�V���Ds;l"�23���x��[8�Hぇmu�߬3�*΀���$͉���%7Nj|c�6���hl�=����
9�Ѓ{c%�e��D�&���4��}���T\P�l��U��Z�Zbֈ��K�{��"W�C�b�O��g��['~�T��.�T#v�%�����
�7����2�;���:���Ԏ��ڤ�)�C�!^��]��Or �C��t�>�g�(�}-4k'�M�h�a�~WD�{�V(o�`Y�9��%�ϳU�$HET�V
8��򏠯Wb��/�g5Z:XS稳Қ������s�pqfl}5�<��i�=z$�1Ze`綡��}2�4�n+	�ࡠ=N��)t<��o8���i�z��Җ^�����6�-��|��52�R�#e ��t�q�>��r����)A��܂�[>R"ED�]�L���}Tǥ�7<�D���D��˲��P},$��,̖�<�Ò�%k&�R	��!T�uȦ&5� ��9��S�[�B�u�]^�D��ycȱ����'7�>ь���sB�&&}��2���p �W�D`��~-h�J��#��z� �-S��\�L��u�� ��6�M)���lQ6��*t��Q�PEfm���(״C��H>tP��6ɖo�)8��3�ɏ1/�F��i�#J��-!zr�9Ю�I����[8��0Et�V�S�CO(���-x��-T(��v�E��e������E�&CX�p��E��~�w�`���˲�JGx��%�TY�|��*]��'4+V�k+�=�" >$+),_���ނZ�
�ĦV+��;91p�,�f0�Q�/?�3�&<:����|!y�'�����en(�����$����Łf�uɌ:z�az�e$o�_�Hm�X�&��o\��y��/�r���C��j��ͼ$v���(8UVS7����{$.x��c-y]a�h��P��jK� �M���Dx�QT��:햆�oZ���A��i��0����:�_��_0��5��2��يn]���������N`=,ݷ̳Oҵ;�f�u�X����GW�X9��.���i��k��oxw��a����[��4H❵��Ĳ�<2s�[wQU7
��|�c�9���8_�1�[#��c�iJ�0j����dT:.N�;�Jlo�\+׎z�1��~Y4�#���혪����!؈�{��\��R洺�S�N�'��%]������2K}�'d-��G�L��?ٱc47�~Z�:������G5�.Dk_���1F,^���1���Ɵ
irϻ�B��ߠb`)��%���(`+5d�S�"E0���ɉ��{sR�L�h�D'��#Є/M>4E�I��$�'�t=X�Q�5�J��Pͱq��#�W�wt��,T��&�#�dGs������3�Jơj��a
P�pdb4;�׸Ǵ㕉hx"Q~2}�*�#�h{jYʎ����T�l9��`������Z���~nNwjo1��pLn���o�N������y�m�V��F��3>.�fٿ�b�����E�>Ef�3�26�����bo���鵙og�~���M������cߗ��e3Fh��f�����s
��#lB�gY,M/��9)��>'k�������}\k[ty^S�o�UV>j5¦68��z�lV�?���?�v�e���+z�-B���N�ҹ���1���6�D"��]��� �C���	� �K?�����W(��zUY�u��Ħ��_m���:���������?O�g��r��$�̝Y�)��&��ejs\3���J�C�׵�I-"M��Ri��5�yA��%+:��<3S�7c�C�5l"�Sn�S$D?O*�T�,���K*�Vϑ�t$Rꉲ��[e<^�d�|>�kc�A|��c|8eXN����~���ǤP�Ц����!v_�#(c�d��=y�إ��"�ᔌ�ͱ� (֮�)����������Y��@��Í!���+�ԉ�A�}��DK��+6>�V�H:�cçG��D�pA������b�%T�������^EW������@�&�@�B��2U^��B�b�,�x�Y� 8(ע�	�$��x������tP�"����WU49��6'E�vz��C:De ��5E}1
��q��a]�v��UaPҩ�Y*�����1Hj���dsh*��o9� U£�T���cwсXpf��d�o�Ì����a�c ��W���S�|�ͪU�rQ8W�:&ϓn���!Ed�W��RϹ����?�a�}�16�PE�m�w����MSCc)�e�X��y���M���$��N�>D��c�G���='��ń喣���;Cѯ�v70�jE�z��/�i����� ���\^]�r�I���z�3�ٜ<�c)�I�����|o#��ӌ#�({m�p���q��e������J!�J�r��ZF�Hs�Q�����HA�pv�7��BD�A^����j~e��\�-�F�Ŧ������T�����C],B�:84�3��d�M���wh����k#�"&*J㒲"ʘ��e>V~H�ەz!�<Q�}�Iw��֩wR]M�ې˼׸'}$cʑ��&u�a��v�'��
}n�G,Ǿ�P�V��k"Ǻ=��E�R�����]8�����B?���#N�7Qƺ��^/���@^ʈ�{n7u���N��Y���G!��Ҧ������s��!GS��>`J.�t@��'(�6Y�`��L����~�NiA�-T�&��ϓQ1�Z�/4���!���k\�v���Y��'Ea� �U���"Y [�\�a���y[t&MtkU*qb��azƁY
�F��i�ZEε)�,���+/d�l4N�쬺� �"����BQ��"�2�?F��PO��7��5�ƤWg�a'���.0�+q.�N�"+뷹z�C�_t�w_�_��'-���S�:|L^�r~�i�i+��Ɵ�i��;��#j4tc�7ԩ��Ӵ(�i5���O���>�<F���Єgp��(���p�bSݳ�}m�� Lg�bݘr�!u�U�4o/\�c�{�bnk!�3q�Jj�Y#����l|�CzvwֈITqOy&�ʯ��[�"e��:Y3O��ʄ�7�W�]�)���>L��Em�p?$�x�i�+�F��������J��p�{�	ydG��G��Gmג�vo1���/1�!p�y.l;Q%����N��{H��� ���x:)V�O/e����;?م�^_jp�L�v���C")?��bd֜��O�������ZT񪒜�E�rR�2��l��NT8��	�XrFq�9��ӬY�Y�ؠ���o��N733{�
ܡ���{�]�+��0]@�zF�c�����.{sB�Ց�*꺖��-C�D���K�d���,a�*�"����H��i�6�-��{i�������e}1�������"��;�^N^�<N��(%�*<��/c���.\���1�`5��f��5�J-�n�ٻ�wH����j�[F���c�P������
"�^bf����U����@5��H>��@fOD-2u~/����<����$:@����f�#�&��+f���OPr���{0��6��q�]>?*^�|{�ǐ	�]�����~?�WW67��b���Kn8�w�B��*V�@`(�Z��MM��J��Rs]��R�j�1�Bt<�l�I��qc�U1�q�E�yX����}̓J@��r���r$�<��]R�ܵ�Z�+�������޴3~|��g�R���Tr��d�`[���L�+V��c�:3%���*�!��0M?���"Gk_��w���Zz�,�g���t3�����b�cPMW���XsK�Ţ!Z<���u��y�Y�J��Pp!������r�>MIƺ"8(Z�D>��`�d~��,V�c	���K�Q0C���,zV���'�#JL��庰m
'�<�
����h�^V���C	5dg������;x�[��@�| λ\����xd�B����]��^iVW8�yŀ)?��d\?V{/��"nt�*�n͎ >�G|>%�q^H&�{9eT��:�g�����ڛY�jF)��X�Sp�i��p7?�˹Jlp�9mL�F܇�*�vWzB�<���o�벶��Vl�!8�\�}Ԁ���Q���m�{�@V�DK��v���w|m�3��,8���ݬdR�q�{�=NgO�s�Upw�r��4DI��7N�\#Y��w�Z=?
N\I�J����9@�F&V��sw�K�Y��t�d��~;8�RQ�1#�ao�g��#�="D0vD�7��&�����}Cx�$��i�O�#��OA�|NE*6�t�k5P��]�������z�B�@�7���o�w�&v�fb�p's��Ry�y՜�;���U&U^>h�O}������ψ��
��=�=��z����V����c.JZ��0G:Z�Tr�q���	P�f������m>�l����g�vM��c
��Ib��((�9yɾV��!��^���@�7ў��?gHe\�Ux(R�RjG/I
x��z�
�9*���4�)�J6��0	���i"��/��#�$1w,Q�*{��Գ�7n܊��jAF��us�6B���3�`�U�������w���L����8�./�B��C�J���D�I�dJ���NyS��{��ۣ:;���\Ȱ�P��pP x�X�QO��t�3�kl綯��u�Z���Fj
X�(��7~e�4�KN����`��Pt$����<��W�V�.�]���V����B��.�#c��vd�4 �d.�q��w.稸(Z�jv��	S���`�k�mj��T��b=�u�� �MÙ�U�p�Fؓކ��o34�2�o��G�"�#'-�^���r
U�Ju��m���#��J�PW��� �Uh���9�#r�������4�B�	k|�s7�����M�S����C~�Y���sN�5Қz����w�� �M�G��.�_�v)U����@L�x��̱��u���Dx�.��鮽����S@z�I Q���5C&�9��v��qג��I�7�O��O�������-��}��:��/_bjK�Sl�L�R���tZ� ��?2�t�VO"������w�����S�L�P�Ͳ��T�<S���T�i��ڝ�2��>�g�4"�u��,�� ƓF�#��Y ����E��ʻ��N�	b�j���N��A��9N6ṇR�s�`dL�����X�p��Nr�3Y������MLI�=�DCh4�a��d2S�3�3:d0n�^y[��q��~��*����ͤ^��*mv�j�.qН%��n�ވ��f+���Q��l|����ۄ1K>��u:C��uL	��f�丯��ˎ�0����oT�Xe�Ȗ�#]�����^w1�7��𘶑�	و��HNf]#m3t"��H t�aq�(x��$n�穣H��%��Ȏ1&%|�Ú&qHG����*�wBb��FI���*�^)�����I8����u�� �'�a�3��+}�h���c� ���������#T��=�B$b� �t��aaU��Hڌ�d_A�bԨ�O�.ň��� sz������'j�����S��+(�
�Ԏ+Wv��ƚ'�6~�����_�U|V��zAS<�4/��ˤ	�/�~H�V���n+I�F�"��ٌh�#RL �����x���e����1{-$�zʈ�m�e�&=u
RA�����=�g �;ژ5j3�xoEn�6�&R�>݂���SBC�����ri8��R�R�t�N� 0|)A�8�CGe���� �_���TL}�b��6^;L��_uX7S�����e�E�W1#ؐ�%k�}��x���B����*����D��fv��~���Po�Z������7PE=�*��Fz��\z�8���k�L\��J�FV�����|<�gf%�c��)�j�z���w�xM�OV�ۊ�xi�\�7��������[��Xm��F�F�~��9�&6wy����ud�^񬶇�ӥ���Fno������8�C =Ѝ)jC��N@���K4=(���ļY�H�qe=�|Bn�ߥ�П��ų���뾍�Ϭ��O��݊5�����1�|���u���,���>�Z>9��o�X�R3��wĤ���[�6�\�3<n�vP�o�m+R�
�����8�@w�7_'A��T�I$&1u�y.Z�$N��m�4�M�E�=7�n��bpn�J���jΝ?�7��������A��NNpIc�%����'x�+�E#U��e5`��E��"q{�R�(Q�����T��B���/�1�������i'Hk|�ݜ�4�7M
Sޫ�t���Ҹ��>HmҌ��cT�>�ѷ-DC��<������£S���T\�D{	^��CcJ����5V�~�����N.�cR�B����вM梡G+<f�
i�ёn7�9X���\��C��o�̾�q]5���D�zǃ��֯+�J�N��P�m�MK�4J�$l�ƩTRrq_��g��O���E��l,�W/YhY��r)ߪݩ)o�J�9,ȭ�c,OO�;�B��Id3�[d�:�l���
�;"��|F��P�}«����������C�SB2�d�I��.ָ{��M��%���z���a���A���gTك֖�)�>�_F1��8+{E��u�]'��J)BGV��:4s�k
TNS�QS'���ǟ�]��F����n�󏅠�eTJ�1cУ������[_�6c�4�|�ҏ.�Xd�h�	�oN�!���h#6S��p*��'�e����x�4+@֪�I�ö&9�J��|I���a�!T�ܖ� ~�7�uݕT���T�D	�RѼ�(�!��T�A��	��ɭVg|1At؛%(�ץ����<W�gW_6I�Ay���HVG,d~�쳠�����YV-��|���	v}M����S/#*v**�#@��Φ�)2�K�f��L}�OVh����^�7OA�~rY�)�IO�7�gق�Jt"0a)��r��QPF���El�9��X�43���Ӏ����׈6���	Ĺ27�v�?t8f޲!�u��L����7��x!L��`���G��#�*�}MQ|�e�nY�֛q~p̶]����܋��c�z��pb��`�����_3���V�4�A.�t��?�*�1���l����:M7�v@ޥ�J�Z5lnͨ�Ah���y���ddҥ�B��6�J#�9to�ya-*��A}��T�e��v8^KD뚋MZX�ڔ�ǀ*K?��o'Ѡ�����)��a-��ƵG���׹�|�6�(�]B��7z�Ya�"�+��2}�x1"T�Ą%_�R�O1]nx��s�vL1٧;�f��'s�_l)�92��S	e	��r�cZ�bj ,�O�����ױBaN�"!rĹ�,�ss}���Ŋgˠ���?�j���B���+U�n��9���jPYq�ɀ�{��X��rv̉�1��i+~���S�(��9'�<�#g&��ߦR�I9�^>띛Ex�tX^^S��>=	h�s,�x@i�qں�~P}O=ER��>�,2����гNA$�R���/s5C��l����q��h}n�#�!�/�aGҁ�}��}wS��(��!�Z�*p4��Y��ߝ�`� P�/r���#}�!^����U�R�[�Yc�C ��0����46d�"��k�6�	s����n�	����Y�,<� -�nhw��E�����C7�e�W���L Dx�C�>n���7���ధ\~�'� �S-&�q��Iw�ݻ=(\��oe�����i��	tz��ʤ.��鹶RGR��I��x��;�n{�t'mt��몧V1��h3)����{V&�,ϚVQ��E�	�dH��Lӵ�K^I���@ #���d+6����k��Ѹq{_���)
��oy-�W[�AVq�4�b�9`vk�$����dzA&�T�1�bu�c�uo1' ]ˍ����&�ɪ\#����Un׷�\ �2��-�D ���z��a�}�H�f��h,B1�'�,Ϥ�+�B��r,�����P���S9���\-}ʜ�Ӗ��3���k��l���-�rJ�dB(oy�,i�W���i�k�hO��8<{t�G� ���=nڶhC?J�l~ n��$#�J�lB��	�}D������X�H4�x
(WX,�a�ĶbB���\h��c&i�"�Jp�ȯT9��\���3�k$�<�1^�|�7���͞�KA2�(�q`���ך"���0�h�x�U,v��mL�>�ξ�ÿ��'�����.����	?h����tC#>}]�8H/|Y	�T�}�HU%��w�r`Ū��Q={�����g���Yj���Ӑ��de���~������d6��f�{�`������qY��"�潢h���:���4i\�Y��A���"�n�ؽ;ؼ[��XI�K�� MM�i�e ��m�I�7��rN���t��Ol?5��
��R���O���d��#`?������DU�����5t�W�D�@>U�cY}��a����c~@������c9L���!u�ե�U��ǂ����r����%����z,�B/Н��k�V7F}���<��њ?��r�0���⾈���;�(f�����S%@r���%��}���f�h������U�A����&+���Ϳ$R�8o�*��l=���}�?�3D�蘿O��΂���씉�x'���b��)38Vy�Ff��k�������G��9(�&��iề}FTw��$�E��'o#�t�
�av\��C�𖈬f7o:Ty�Ն�KK?���:JЃg���8I H��<�LRN	�*?ώ��4s�[��I�0Sf:B=~{���,=��w���
 �kz�N�,E
� ����>��E��\�Ӂ�jI5�<82��*%��{5^՘�y�1Ȱ�L�	_Q�x�(e{v�Q>���%KJ��x�����;�Lv�6PO �굢pM�t���5i%����g���]�h�]�U�o�5��r6�ۥ��f�� <|<w1p�hb�v�k�.�f"���lj_#at���a?��1e.�9
!u-����yzh�MD{p�p��][��n�ndT�آ6�d�s i���a���8`���ן^c��;H�g��c2�I?��Z��&R}�3�T���E,s��_�GZ�B��+���PE��������d��`�5ؔsPb��D_z�XɚaJ/����)�٢�^�hLԗ����+X���p0��ZsJ �Xث*�fa4��>�6��/PUH�mNB��uD,��,H��Q�|��E��)c��IUt�0w#x��Z��h��f��Ιmfz�����cbJ@\4 �S��_�����Lo%�aiW1=VI6S=֑AҴ�qa7��;I���U�I��@r�p�[��P�0�����3��F�ˢu��|���ȭ0)Oi��ܒ��w�d�DЖdFP����
䄟_�~�n�[�(��tH���u:�J��_A��ĝ(�VP���g�'lJ����/�J���}���P�22kQD���ȯ�
]Ԟ��_���j=���4nzCE"���?f��I�d�ɿ��S0k�V0
|�xd��x����dtg���{h\�fE��sGZn#���0O�V#�%Fg�����`VlC���cC�����s��8i�X��:4�ο��!������HG2�nG��ǭ��>�5l�N�2��h��G6¯�(��*!��?���z��rU@�����}��B��&��J-ȝ�x<|'��P����ZW2@�%P�J�k�ߙo)��$#GJ.����Ɗ�����"��W���h������>D���NxZ����G��f��'&|G��_����/��-��rņ"���:��vy�Y�
qQڠ0�� ��~F�I� ���F�eG����j��-R��P�,)Q�5
�j�^�;&���%���M�;E����(��f�G�T,<8����2�	��J�6�u&䦄�L��e��=�#��ASTO�j���B7�;FO�j�Z�y����߶C�u�9���̎t����
�9KhB��{8�]�mh�*p ���A��A���'�?}�I:p�]�6��p���W�X��	����זo;z�i�`��bCk.5��cl5s�).>�ZГ\����D��T�?������z1F!�R���x1�x��
_�.a w�Ok�
B�Q(	���3�B
�F�rj�i���hM�2�V מ���t��e��@G���I����M�+�K6�Y%zO�� vƘ]�Sy�D�_�;����/8�É�|@ă��.��EiP�_�x���Y�\���C��x�-�-�5�\3��R?�N�fص����c8309���u��[��t�vyj��z�]\��6[��~�˰Tr$��{�u'@}	�89N��ԝ�֤@���2�����:�8Ը�׉5����P�V����{;�[�A	M5�x�m_�n����"�p�V�l}1�X	o)FE�Ī�-���;�I@��͵m�E��E6��p��V�P�@vM6'jU�=�L�Q�zK��̥�{��L��U�:F^/e����e=q�_e
���G,ק��Y�(c�oI�R�� 7�!�+@�6�� op�N[c����{M�I�$:�	!D��m��wY7������0�t�I/�%� �a���)M��z�,>_XE3�5�΃-�ί�u�ַ�[�!�a��>#;�N����uA�e�&�.w���P� �U�@
�����at����7�1"[�Y�����c'�"��v_�0i��5;�%�/�&]~����֥��h��߻�1J����
d2|/=e��;�����x�'Q�C�2
|G��o�l�a�M���W9 R��^�@��V���84@�P��;m;΍�a�o�]��T�	���T����@��-���#�C���5-&��u��[-�`a��=H��0��|)��gW ��|�/�
6,N��{sn����uú�<r��/2u� ���K��d�m�b�?�9e�h*�{/_��T)L�8T�>�.*dۙg�`[R����I4\II�ޥc�?��(Nj�B]߳�I�����Z�N%�BD�d�	��Y=Bq�ֶ�g�0Sc�q����y
ynQ�Klw#���@��[t�g����+$�|C����-U*������N��6�o��ù�]�rˌ0����{���~�L�0�;=�
g%
��wd�_�q�/lK� �q�D����*��O���Ŷ��Jq�_`�����5��UpVЇkfM���t1��l�\�SE�<*i�rjK*az{D�_�P&�%|u��	�!Jcq���"=ժ6�M���u�b��AȤƣ�@;���{��j0�:�⻅dM6>��Z�i����ɠ�=���p����v�z���ÑW�G�!�=��V:�@I�i�>�18�)�������s|���b̉�Q� �p2��}`�\�I]��0����z��h_��v!ޭ�E�x�`ޅ�G�F�����F���F2���x�C��PP��O1�J�^�ێ�\���tK�&�&P��e���Ț��ߑ����_#Fk����v�71�yhmT��j�4TNq��o{�v}�*��Й^�R-McHgWV��2��S����_1���BKrF��A�}�lQrtnc}!��C�3P2�<��"��1�$����hmKu���XXU9�-�A��Г��T�t��7?�ؙ/-����0f�$-�!�UB��[Qa���B^,�=
��5�l�"ȏ��rK���!}�rJ��˓W����V�'��w<��TZݸ&D�O�ӭ�6�}ƶV�����R,�`�C:�4fh4�x$ܳ(�TJ�_��*�t�3�6�'Rz�����QF��b3D�.KfY��[^���'ҫ�X��t4;�츒+��>ök�$|�,Pb{����dN�h-� 8=��va�5�Lz�����������IbcKWE�e�Q��1�<�_J���N� ���I@������3�������!/+��_ϊl��*�ܰ��/�s����v��ULk-���5Ƭ+=�� #ª�����AX��ch ى�9ǲ+�: -�8`�1�e#ؒ�e� mm2����ǽ�-�S�N�0v���b�ldnp{&��w��P�ª,
�΂�n�����+��J`�Y=���5��?��x�$OvCʂ��6�ѯ�1I{M�����Qca��-�.�H[��f���� �yG��\Ö:��']�
�(z#cȽ��y9=�%�e0��]P͕�-��qm���&=;��7}~w�^� \^�����!���B=�QA!��ʋ�Pʯ����g�3*��8@����Bm$�F
z�L:8E��+m!��L���E���������Vǝ9�X��m���ƥ�݈� ��/����\U���[nޫ�`k�.��.H�Z��4~7�/z#d�0q�\2?ɾ��$hZzwC�S+؟����E����t0��#��샏�":a̡X ?��oM6��^M�%�ʅ~��f{~WQVޭJ��Ci�W.� �RxP��W���:DV���ڪd�*�󞵩B�p����\��l{�j7c�����Yr��Ƃ�s����_(l/�����\Ƃ �E�*` �~���T<���ns"���,�]�3��
����k�R�]Oɘ��an�(��R��h�+A������x���*R}���f������_6����
nf�?G:?�n!ܴ�2�7��̃-5�k����2Z�p�,���VC���c�R��	�����;���G�%/Y�� d7���$|'}甎W
}����z�����!*�:*��詎o.��3'(�F��Ԁ��t;L7���G����b�Y�1����͑Zf��dF���<���.�uS�I㫝��z��"u�"�x�v����\Bv�a��x���J�94����.�mh�
B�To�T��x(.n�����:��C^���m�e>ت���z��6�F����br�v,���}���eBd
u�
P�Z3֕a//(l'�T��ոt����J	����u1r��7t�3)Ũ.|-�=�����&�8��-CM��Ә����/�ޣ�dekc�Ӡk.E���A���Ml*��ّ|8қ�0�q�-�j�L�u���𭝠�#,��p�xt~3>%����-ژ����f�,����(���H
B�d8��7��Z�(��# =x (�� YN���pM���E�D��z,WG���5�������8�|���2�b3]�_�l�o�q��=j8FM�_,Qc(��Iat�-�a���0���[A����Vǂ?D�����P%��|"��`�gZ�k,(:)v9��$p{֕�I����Ѻ]��k9�:����d������ `�2ʣ���-�8��lʸЯ��I�{7!�������RR6	ODR�}Nm�\%��|����>��T*�'�lZ7�|� ��:��������v;�Xdh��*i3�t�.�~�C�a�m��)|h�}'˺��6��<�vo���G%�&[�h;�#�G��D� :wĦ������M��@�Oa�����DI�ϱ�z�M+�v��F�6X��~&~�(�*Zf�L�!^#u���B���>;���zF�3XS�QV��� y�����,���;+
hS�i2tB)@M>�c�z��ʥW.>뉶�����=�6������{)�Y�Ш�^�&
��<Y���jt,��¸��J|�U��˽P�)b�n4�`�_E���\��U�����9��t�|�Q9.V�f�} ��a�&~V"q���e�`������ɆoD�� ��u
��*�xQ��*r�L�/m��uD���ǧ�-��l<�����KE���>��f��>�Z��(]At놤Y���5×�k�׮�'������2I��Z�y�����x��o�LG�Rf���'��jh9�-ٽ��]���W��.:��MPX_������)��R� ���d����D���g^��^3���-��%�	�:�M�^G��7&��sQ�G �sw��Q�d5�l��#~="�[�`U�p������O��=$�g2徸FC�<�d�^���V^^w��,����4�r૯����$�pW��I�!k4�h�d�w[f&�t�h �&�_�?�4sJ�L����>��وdޝ����Q�ò�?�w�㠛�2�5fs�����RH+U����}M~��e	�'�?���g��`�05旝U_�ř� {O���å�V,�D�z�B�����b�ķ����ˍk���Bb`���jx �t#����X�Ԋ��l+�̰KDr`w,�l����3j�����-����?[w:� Iz'eE,,�g�N��Q��,�J��O�ɩń�N}�
�4pV���A\ߝ:���H���Up�_���,9��W� E@�0D$���2�U����|�g���?���e�R�16�%����_|���;-�L�>�u��T�̅}g�U�����Zx"HD�
o�,�Tu)�������U���	��[���8y膒G®]�rᏨ�:��|f�[s	 9���ړ	!�i�����}�Ek�V�^��	P'R�g<�j�k����$�A&@>�̇�cz/v� 8���6q��5A@��#�V���n�z	�qm���%L��X�]
�^�5��� P�9�*����=U�:Dr}U}��YR���%�MH�O�#KĻ�\A+2�e�U5�D�P{�f�a��ђ؏T�ՠ,���O�
�$,��c�͎��ef���L6���k�2�|x�G����,=�i鸁���2�F�S�i�M�^�|��%au����.%R#Z���7�`|x����ʐZP�ų:7G����_{�uևVǺ� fv�â��J��wΑ�(l����� ��H�nq�r�gm��\߀��'J�N��D�^��sg}�ܴ�z�8�F6z՘�%��Nz0���v�R`�Z�]��b5Q4���م�@�;~*on(M�9�B<k���n��N�G2�E�%�ţ�w�σ0�g�9��WEw�p�������pp��8J3�� ��X�}W��_u�Ix�C�|)�GnDл:fGhT��+�~J�Vӆe����[F����էlG;��f��٨�0��W�rִ}�r��5(�P���}�Ҷ�g[3N5n֧P��V�K��֏����Z��֬��w�1�6r�Rp7�n�&�o��6c_����Kt��sV!:���D�j�]����պ��y���Z V���ad�6��#�u��'�K~�'���B��P���������(o�t�m��`��d���K�A|��j<f�>�.��d������-R��0w7�ݷ}��U{AV�'c�Ve��f �u�]�e���\d�����gOC1U�L�LP���=�|��j#O���E:��H�񼝙/L������i�/@��_Sa�a�<�a�{, �r�m�b��1��%�p\`���,"�h}��$�E����<�Bxk	�YM����T�����ӱ���*��{��<^�!���F�[E��m�v��8��Y=)5+x9�j�]��������ζ�P��S���f�pǍ
���*Ӓ}���	j�E%�±9�����U����	�k#�%�ΙZe�ep[�RT�U�i	���+_����$[�N=���WͰ�v�!�f�L�w�~�������h�,T�P%��K=3���[a_�W'j�����dn?�K��ڤ�v�A��X;�Xq�\���Ԑ�褧zm�ʠԼ��y,��#.�U��t=� z��_y��Qt�\%�B�׬�i0_)�楥�FǴ�g���=}g�I��grS7��cn��F*,<�&�;��EU�t:{�@�gF+�4ǟ�,�K��1Gd
[�Պ�R?컃7��#T�$���f���W�ؑmk�b���,�!�k��ӕ+}um�i�o�_�5l(�|@�\uD�����Z�5Iݐ�'U)���zJ�Q��Ik�1�GP���LnǪ����i��~�(���H��$&g�
�dg!Lf~���xUj��F����x��iQ�n��FƦ����̆�ܾ�(�O�܆�+1��J�l��WJQX�J^���ʃƾ�mKH�K�����5����W���+�P1���F�O���A�h��{��&�O군�	_:�n׿�h�e�|��H����ȑ�j����6
�*��Y&i�y4Կ<u�֭�]t�Է���L+W��� <�cg����׋U�g���='��4�x�<�jiv3�n�TZ�ގU�"��%� ��s�	�_q}=9�Ƿ�f����,7�#��<)X���;$ȅJ��.�cH7����q;ep⍤�	b��3�TD��? ���E�����o]���S��o���ja�m�6^<���N�;�Qv��c�Y7|����g�xc@����٩�$��FrMɕ���c��E���w�<=yߴj͋�ը�h�Z�:����5���Z�@�:��.��$��9����.�/�*����E��Y���1#�>�R)Z�a�4+�]adk�j0�Kl�~\���������K�F
�n�B�5=��r�L���
-�4�P�y��n	�O8�kEs> \��:���N����9qQ�5=UZ�*Eo�Ʉk�[��Z��׻@�u�+Az���`���A)1NY�t�5�km�72��.��(?�[c�����*�$���낯��U�*�bp#*�/&��S���",���59jP���S���t��=)��9@�r����ǉ����[�j���(�S�>M��S��^ �!��q�2��K�n�"��`�#�dj�d�֍P�!̪�\����ep�����[z��&ʄ�Mxs��������Œ���ƺ�ѹg�
A�fw�c-<�u���a���%��?�	lѲ��R�?�h�㝌I�3lX슃 ���ȵ$�oc�����O�:�"́<�Y&��i�y�m�9�ɤ!�񧼂��c)�+D�nr4�"��n��a�Ԙ�B��\BRcW]�q�O��Vl��I;+�o�F�#��|��m�g�	(��u٢���z�}�rÈsw��; I=)�眾?�ar���s�K��1�q.u��ʤ�c��B3�R��q�j�+����4�NP[	�Z���bJ���i������Tm��Y����X�znʼ�]��M��&�/�ߩ2(�v];w����i������$LYDØ����p��j{"�O�/L;K`a�r#oQÃv��}��*̫�nP�-�&yl�7���*�X���O��ʌ��Ot��}wM�cb�u7�7�1����A����SN� ['b��v���N�0 �e����6��/��:�ﮗ!�c�#9��i���I[��j'��AŚ���p^�M�������#�����Tc6j�q/�$��/�`�n�c�)�WM�fc�I�8��f�~Y��`LغJ��cir�w���RSs��_����[���ߧ�L ]�od*G>��E�!��;��ܐ�v���ځ�b�Ŧ5��Fnщ��W톳3�N�0y+�uav��%����j���?ϙRΫ�Wȟ|��Q8�^��X���k~���.>M�e�^�@�y$Q����¯��4��
{��S�W�$�1E���=F.��ʹ��s=�p����arDz�W����x�����RI�=��w�6��p����:6��X��)�f'��t�R��`o�=�X�W��2��K�p�o[��S��5/����|v�WW�@�&�L��Լ	��^�C��˭�9�6:�Q��D��5$�"��ɡdf&gH���Hj��T�B��+ Ǧ/�3n�ž��2�Z(���U�M�L����P�@��g[O���CyȬ�Im:qȊ_G��>�K��g���БҎ��q��pa�`��1S�Z�S��>��;�?������V�׾�RH��MƿGV� M�d����V�8��1l<�L��`���ѐ0��rT�}o6�s�m�
��<�h�?���۱�r����(g� p�����2��zۯE,�+�gڋw�!�������Ԗ������77rd83=������P��@����u���Qy�;Y���4��nִtFtc0�GdCY��
M��?}S��K5R�!a������B�D��X���D�Qv&)���@�_����,r��e�M�2�IH���%r�ʰ̓�s	�����YЀ��뭙�,߇:�Tق�m��Ѵ�v��G�r����f7
O��΂��/i#.8\ ���a��a]'�ƞĝL�&�;�7����q��G����R�)bXxC_�|�Xn�t��UA��3�����{n�}&���6��*��}��x5�i�u����r�����&���L��5�m��lL���bM���Tq�V-T{,�O����hm%��<*�и��^|NJ��#�&�<��D��%N�x���#�WQ/|#tUS�pvm.Ofsm��6��'�%S�3�/��̞�>0�)��~2����y��Fό�<>ە�y9��j��g�$x�Tܯ �����k �xo��tLd��]��E����C����5L�����J*����cU+������S���6t�Z�wM� ';-^{WÖr���U��I`-3.�!��fC$-eÉM���N���1������YH�����,A]�3��F�O��L�`1�?������Sq�sZ��!1�k�G�1�vTBG��4��=S�\�p��7��Ǣ�kõC�{�@9%�<=��)��z�+ԇ��vv�J��0��&'��s0*�P�	�9�D7��c�X�?�:�-2�_���k�����çv�0(!a�a�P�"<���A��0��'7&�!�-,�huDC��	e�H��m>��5h�h0���7����,�_Rn(�ޥ++�;`Z�/���(�=i!��ǥ0���?K�Խ@C��?Ǒ�0�s�g���$	0	-�yX��`¡!�� O�D���q�.���2h([{7��Y��g�����\9�1U5�FR�{h��bD��6�6�۪���ؗ��e]-sh�Pؒp&�:N�P?�����ئ��X��m��)Z�h��E8,�5�����b�k{���,G��6�����6b���̺�^vr>���Ҍc�
��8I@Sys~Q�1�����r<;�|2��Z���݌IgUj􏉭��-�c���Q�vK|˗��{t����@XR�w3�>6
�^�9��b�L?�kS�ՆY)I�}���6!Fm#�����]1f���J8�� D�O�w��@_߷T�����׉ƈ&����Lb����;\�!����t0�'�X�����b���̾�����
�q�x�p���[ ����PA�JPlv�P�AU�"���H�6�rI�\�x� z6�����8��T$�[e��W�@�W����ŧ�l�8����ܖȿEQ�Ϋ܂�f��x��LcÂODO|ی���Ia�#P���լ��OhD:��+�γ����7=w)�Ұ�~}��"봬u�����e����}μt��)�� [��������U����UX"���WƖ�G��=�@�=܌ж��@M'LnW�����Ĝ���W �Y��-��g~��a� ��$R���sr�v�!��K4�G6��/D��O.up͏����Y��G�����\c{Ǔ@9D�{�g��YO�$-d�!B�r��my��2��Lf���q���h���`�&A)��J��=�ڗ���>[D皃��Z��։eK������fat=w�k�qo�Gy)�g�'|&Hy>b`=!P�J���������j��:�^_��F�h{B���١&�Z,��Bx�h��<LL���"J�M@I�\���6g� ��6�.a?�$��-k�����M����H~o� �dm������B�T�ΏQ��I�3�^p�SO�΃��x����X˄�P�?�D8����{�pRT�Ƃ��v�ԅz5�-[��Fᮝ�Br���pU��#b�|�Cd^��hЌ�eDdr����7M�,��=�X]���Ԡ̱����G�*�F��H�������%#&��e�p���b��bt�k�0��'�Hg����U�+�G��� B`���Z-��C�?�.��Ή�5g�gQ��ϟ�>$P3�O4�G��b�����5{�@)��R��Na|JR���Ol��3ǸV~�������F6����Iĝk��B�߃�@z�^LN��7�2�b���e����JQ��d��w��J9D��\�J��Ga=��y9��0� gM�a��ov��+3���3�j�;�1���าå�)`�ej���ҙ�(=�+�I���!���-R�,��o�,?
�ID��q}싎�D �C��u�Òl��J���0_2�q�c�=R�O�VZ�jZgs_mB��' orWfق�mܕ��p�]���w��9`����'�:�'#��(��|�P����K�M\+���-o�mlX���F2����]�J������'YD�)��Qp��'���O:�$ �<c�_�=R�{R����௚ܲ^H&�Z�l[;��Foc\�\�ZfM�ٯ���g�C��ZPs�N��&��l�L�� El ����L����W��+u�f�QuLZ����59�Ve�i�Lh��j�GX�8�_��'����E���p�	�{�u='{���m���|9�(C�^��T����^��L��8�b'��g��3<�h|S�r�ʞgt�!��sd��H���s�'Qnm5�a�Q�>
Np��m �l���<J��?���@���C��]�8���}��:A54;CF�?�ɢ ��j���FЧ}������@0Y:��b��p�Y왥���˧8ƕ�kJ��{�Hc�g�52�u�}V��.
tl��0(޷/�Hl���-Ig�&Ɉ��D��J?� #Yȓ����IuJf;9��H�UpvE��z�Z֑���aRW�/� �}�N@vO�%�����8��v�f���)A�?%��	�*���alUC�7�3�uMƿ�:IU#������UR�oEb:S��D��5{�\H�V~� )�[ˤ�l�+�*�//{9&�8��#h9�%��Ĺ�&
�MSXӂ��ʐp����cj��]Y�����lW�,�a�������o��g�o� ě�,o���i��L��Z���8֡��<<</ڭ�#Z�N�氉,�t��X�\����)��n0u��+��^�e�{dc�.��:��,�v62��tEm�D(O�����@�Z�<<��ʐT�ٔ�B;�[畘W�T!kx����#�w�?2ܖ#��s� s�(7�25��9`'fKH��=ss����w��o#J{��E������E/�kX9�� �&�Õ$����Փ*�|S����C*��+Fԏx�_a����[S�	�B�B2dVғ��9�y�� ;�i���ʤ/+nH7
i�@{��rD�4����8�0G�]����5;$'e*�������S���ޑ���S�3����ŷ�Jf�}�qLg���"�6�^���ʛ	�̾z],������E�d��#?�>�<%�����x��<���Nm$��������� �lug�65��<���*�����[u2XKq���� �h��+�+LVٓ�f�8B�._�L_�������d�mgEB��h�b(Ճ����J�DGD���l�^���u�	{.4S��2�5�������ۃK��$Є:e��Mml�m̂%(Pp���}�XL�HJ(��m����z}.o.H���k��Շd7�!4�!��)29�I@h}7��������>�]��a�L,�{�|�7W{�c�����h�!\�RT�5�⤔�G����_�4�H�� ��)���1&�sH+�hW�elY��6��&��m=wn��j���Q�iD"�p����Qf�+P�ک_�z0�G�wD��P�_kWjaw�F��Kŵ;��J�?�}DTt&ڌ-$�lʀ�	���^/0YrOM��pPd��Y�ш�(�4֧{�+���8ܑ���K�DP?VhG���yA
�lL�Z�HY��z�C̵��l�(B�)(�����"�Id�c����:лm���WQdw�tո�˘90����jE�������q�&{���w�[��E�|�TI�@����x��u�]��G���AX��m�,}|A���%�c���)���	��d����ٌf�Mk����?��ױ�.�a�f�44ڈ��_)���K�ڻp��6uG�a����=�t��4�A�W�/K��/�={N��� '��m{�ݐE)6T��%�J�x���,i�`:����bJ����*����"s^S��$0����bz2Y����i��@!�j��M񼦟߃7�?I��D�SM�x�:Al���S���Ȇ�11��{�|
�ZK�a����6 S�Ќr��HԾ.�q?��$yj_�OϾ׆�IG!5C�n���
���`����wqWgn>EzΜ\4L��{�ԁ��Hv Ak�0˰�*��8�=p}��G�ǁ�T	�V�R�b�	���NSi�9�m�a�N�>�)���p�'bM���s��/+�K�����<�9)n�!�djQ�z~G�b�;4� 1�����Z�O����P]�❻y}�:����y`#[�Ml����"n��'2�L����|'/��:ذwvg�����cV���+�p#�Hr�gZX M�1���w������w�q��rP��]?�`7��HX@s}�'"���D�^�Y05����0��ll
l��G��f�=��ׂBQ;�O��xqzw�ߓa:�
����2ݬ�GVoyy��N|��D�����c� ����u��fq����L�0��S�/i�	ǻ��։�����c�,G6�z�q4MWe��������_>0�d���qB%�J�x��+�V��=�C��t���?,����i<�a��oZ+��C�	p�6�Gꗂ��=�w<�A��v���R�I����g��"1r�X�۱k�|�R%*�A���~�eN(����(��D��3����D抄k@���Pڂ��=H��������;O�](��ӻҞ�J��n9zVkDA9J�Gx�KxyJIu��GҨ�(7����I7�寰=�$�i�3��A^�!9�F�r�סּ8ԍZ79,���N�X�ѓ�u5Y���{(��� ���x;��83"au����4��"""��$~I-6y�e�-` !��K>�Fb7��������EfF��|T���SǏc'3�񭡷b��A��ҧ^�������:�=B�׈-K�+��[��34>��1���p�,G��q��[����N�����~!�N:�v���6�	�y'�!G�2Xu�T��N���:)ŉڍ����5̪��$�(d�i!���q�s�9*�܆�E��V�99#����_
�t�я����#R�B���v���,H��3��YZw��g_&��fj�X�$�e����cKw��n
C��r��ٕX�b��������b���P��*�O���ο9��bAc_d��m^�N	���_���`��&���X.&�v����À\@�'5���9؋t8G�ng���:P��pxaU��lŖ�ݍ��I|#sy��գ�`��̨�3V�d���{$3&�[@��+���cW+KL��9j���������ʻU*�
�g�Ɠ�p�iI�l�kʉ��:���9�W�����ͳ�;���cگ%��/������n���nX��0n�A
8!������B��=¬4�Yx�tQv5IVyƁ�G	쓶l�7�]�<f�̽����4�
����%1}R�?�	_��j$$)}��:15��# 1�E0[#G��>M�3�G� 7G����k:���e\ᇩg/`�Θɞ�C�\D+�<0��̨X ��VD�n=����4���^t��B�c�n�$N;{��h�'3����;.�*�s��u�أenR�tn[��z2RX�8�l�D���"�Z_I#t1 ,�����\���eĻ¦���Ɵ��a��T�.DǠ*F5thQ'>�ˎ��i�R+չXϏ'V�vIw	l���Gk��c�g���������3J�k�Hȩ_{�:=��TC Ue�\x,��^oK����c8�08&�;,4�p/P- "r8���H|�p��3*��D��L�U��b9�ū_�B(d2$A��g��̋���^3�%1^W!Wǈqh��*@Pa7
6\1��n�����O'Rc�>��v� ���9�k�/nvʑ�8&�?���o�9�9��u������[��%�`�gl��q�����I�+�Gev��F��>��RT�EOT>�U�k����.�2E�+��E���*��ꖼE)���m!>��)3��,;&�d$���=�,��'nXW�P�ﭨ�� |��]�A����WY�3��z�@���h�Dߚ2�-����; ҂��T�軪��-w5�(%ר�>T�IQ<|D� ؁*�t}�`��In-��Y�>�i�2�r��6͢4-:��sLr���@&3�˘�R@��]ޱ��vԳ%{��Y�~��2$�_���/�^��C�y�V�u\d-O\q4�"B�!��[���\=ٱ/#7��y:��{���O�wa
w�<z�Dll�{�	-��z�Ҳ�1���C�e�:g�ȿ�6��i
�Mh2c��sAw�s,;������6}{??a)�*I�/�k�X��Fk�W:?�u�Eo����Pm�E�Q��6R�<2d���9���5��z���6:��},�F���X�j����}tK�ݏm8G���p5PRQ����놈���f7��7NQ�0��H��AćF���ڞ�ب/��[������͹�d<�QP�Y_�X|W�ME1��y�@۲i�u0s��Ĺ�hӘ��?�z�&�N�<>an�,s_���90�P4�÷�sڊ*]�3(�t�-s'�G(�9R��W��&dL��G���_�h��"�6����ge}�kF��d��Е�����i�ST"*r�7�O�i4l�k4�iiJ��3�
��!}�S0��NxkV�<9��+��BUsU�����z�����m�c�A̭l��ٱ��w�W��IAz��ή�����նc�X��z��5e�'��F�K����A0KH{� 0=Ƕ�l���`1���ł�����ö��:�>& ��x9�����b��&A�A�V�Xb+`��h��p$�
qh%���>pG�h^܍9+��0J������Qfc���3����q&ݑ&rIg�x{��9x ���7Z���}���$!<s��d�z�����Vka���74��?�9�k�ldj;�d,�ڗW�-H˷�RV��Z��f��p6����c8R�O6^��
��5��k<�o+8À�Ͷ a��S�1�h��($)�g�k�r�=H�Y2�.b.SZ'D*��������󾖥�~�2��;� e�F�r�� @#�vex����\ �CJ9նT�$��g�����/��;��b��&�	\��mGZ�G�s\�4StPj���%�՚*��g,���Oyc�b�c�\�=F�^^���g���o%�d���I'@v�G8�r��KĄ2�gj�s���NC.���;�}t�B0�}��ʀ�ް�5�A��J|�L���Ɇ���ѷ{���R�X����~��o ��2aa�T��>9(�L���7XunC����q'�
��K��3?���Ds��:�Gi2&���G`�-l30a�5�3�,�=�h�t�����GhIͳ�t�̑#�5�<��*��E7�^-E�$d}���*1���qbN����[):A�1M}N(�d������+B-����Y4��x�Ӱ)H�$1�?Y�6(��+�*����b��+o����p�x�U�mK|���X�� "	���o����OʑU^�	�~�+����.C�ʜ�Aݓ���I' �v��`�)F���YI�v�BQ�zĬ.�K��q�z�n��_;�B�����'
<�$�]'�yb����3$$64G�F>5�!�'�`b�HTx��s��T��|����+Gݫnj����D"�+sw�Q���}��Fdf'�>O�lvW�+��Cͱ�2=���
�N"��׽eT[�h��~{$�����z�> \B�v�2����7��@�&�@	J�]����jJ�����$�eGB�S9��Kl��s�P���m�U}]��vZ��Bg�}J�4*�Z3�$L�c2]PI�s1�io�<FMۧ%�C��d�L����q��E�K6P"��f���}
���j���|�<������`��n�By�(��/�@���Y$a����F8�E(/�a������8��j��4�m�CJu�s]H]=�Ndk�T0(Է[ƨ����}��+Y���o�
�y����(��[�#�zf�>}�; pT.�����@���P�T�$VU��}h��DnYڦ�lP��{t�<���*��0G�L��ևlb�3��ͺ6�]��0�����G
j����+�Twֆ(��E=�n�J��Yc@�Ѡg�L���Y�0�����W��_U�#����,�3�Д����XIP�`6D��o��[-m/cXb�%��K����b�1v b�^�-���@��W+�G�\/}f�.��Ԟ��b��c�s����t *�+��'�`������p+��?Q��"��� �1�e�m8N�;#���۟H���S���:�%�����T�s�X�,Np,�W��{n����k����U��j,��|J���cg�"P��Xh�*�����`���d�"��[]:�a�T ��=���Jg�J=�9p�^E�}��xWi���<2��1�C�Z��c�RfV6B�y�g7�HX-v��9Y�ҙ�M@[��R�-%���p��/��I�+f~�S���-b�&���:���y��~��DY<���M����Y\Z� L̡�w,(i�@�h��Qb���`X;c�� ��s��w1���i��-�c�FȺ����M�z9m�9*K��@B.�áH�����q_������҂��q'��鷳oխ���w�����Y�cCn�	�
ׁ�l�t��5:�'� �q�@�px��~�t��&wh���1����;z��g^$��0��{�v�C�8g��Q����6��+d	M(���[q�jc~�Zi�#�mj 9�M[|�F���4^���ғ�3^�5{�lR����^� n��+���3�% Ъ��_��c�0tS-u�������Ҝ�����{�:t�nx@d4�x����07��ndI\<8���B3oRBJ�	��!� �����ϟnזx�֘7e��f�Gp�_�����,Z���)w*N,v@�,S/P���y��%B�'Ǘ\������i��/�V�hK	�C+��,�;�x���0|�t�)�?���<���t�Y�-v�y�}�Wz�(
n���H���7��G�R��	�60[z�r������޾PK`ւŜA����=Zy�O�7RO3�A���.wń#�lѵ/����	ģ�9�ԯSR���ú�g�?���^ej�ڙ k�B����"*֢u,��9�o � 
���e�:ƧzI��������*(iD�A�coW� wdT���K��b[�`Fk�$^��}9y�9ǫ!G��<1��C{'	F����wA��25J���NBEt��9	�"u��1t1�>4�)�E7#�J:8�+)R�N�NU���dm��;�GwM8�l{ӵ��&��u�^�tT�s� �VS��}u�X(N�nź5c�ًh)�;�鮧�M�r�07�U�q��c\��A�y��a�}��e���.��6{�k�����`���(�۪�,�0R�.��Z`u��c��?��Jm��k;~��'i�����/:� ����l��(&��m�G'-N���w-Є��E>��}J��۪��u�f� �p�Ղ�P*|)!�4��%�5A���& p����Is�c�
���]V�V�I�=z��5������pȅ#�U����O-��]J֍fE'w�ݤʠ�o	�8�l'��~,�p�5�9�d�)h*;)���e7�;�o�U8��]�7z�!�����i�l���m�m�;j�?�
lȴݲ��@�0Y�7��$k{o��އ �",(���~��}�ge~�1��R{�E���"p�ud�����h�v*W��9���9;7���PNE<�-��=r�GH3ԭ�����Pm���HVl�S�p�^��i`�&�r寋?$���h<�Eȃ�ֳ���'�~�ΗY`�8s�E�����|p9� �����G�
��֛�i��]r���)z@�,�E]�$���`P�5�o���:٥mV�L �I>)�2#���m2o�1���=|y�f.�h-
�����*廣T�[p��uqg_���^�+ B�R$2#�a���B��M ���HS��ݖ�����	u��_�E��T�˚X�3 ����7f��Œ6�q�ŀ%ɺ8B)R�`�Q�W���1k���"���e�T�gk�{ѧ]%Vw�k�?�J,}�P)���Ei��x=��'��Pz���7�{�����3؝(Xa7���ONnA&�	�w�K[�%(��(?d|��^,IƝ��7=-��N����w����!!@w��_jt]�F��oC��(��]8�fk`g<�k	���N���Z�Q��tΓ�MWYz��y7��ro����*������RVIR�h�A�Q*�#p����� �~����b���mf�R*���U�-]h9��,5|R�M@�/�)`�)u���s�j�ӱa(��8cuW��T�d�Y������],}�J���㕗<����a�v�'���vC�1NτϚ6�N'�[��Gȵ�Ys �g�K��1r�ľ�ָ\�/�'`�ʞ�`R�qѴJ>��v代��e!i��&<��X����g������9����(�WT$M(�fs)����-��/�s��!o�.�u��4~�CW��`yɓ��Q���y㤛�[��Mwb�+>H�Ů��]��/rQB&�I�R�tH��������m�x5Č1軽���N=G���<��%��d/���B��g��u\�^��R����[J�)2}/T3�vI��A�@߻��L���ot�[Ӓ$���n��d�)��E���)S�:�a�7kf��~�vg���Cal�`y�1�K�U�$0}K�A�d��ô���;���+R�wDF��=�/��=[�ɣ5�����h�d4���_���P�O�lѱ]hS&F���jf��0U':�������0sgQ�*M��h�/?��*��޹�K��K��ܟ�Vgr�x�z?��z��*Q^�V��Qw�e����a}�b���x���c�6�Ձ��X� �����7��p��.��w���JY7�w�g��As����7O��b槪,���4��Ĳ�[�HB�
�**y�}����;9` /���0����:�3�+GK�i����|z��J��[	�����T��b�rN�⚢Y>r4�3�P+֎L��قC�xc��͓ѵ������cX�&�4�#�b&���$��6b� �L�
���o�5���K'Ř[;P�VJ�F<���g���Y��]-!MkL�����a�N�[L0��&%k֛�N69�m��@�ڷc������X�7������B��a��6�����F�@�V
�yk�*�"�SȀE���2���M��-�[�++}�����V5\�5�\)	'	��)�����@2���DVO�8��W�7�\g��i�N&}
�	�Ͽw�����H��u	+��|�����	kSz�q��a���� ���^��\E�e�݈L��x�P~�0��Y2�� 䕁J��� ��a���L˜}�xG�*
R�w�Zc�� �;"$v��sѫ?�.͑B8�!�#eͼ�wު|���v@����OL��]v�j�}~����#��p�4B�%�����f�\��S�:�B@~ԙ���	+[I����L�ڗM��g���)v���"���CJ�&���4R�eFa7�V�2�Z��N�{x��<�)hK���W*S?9d!�xo�Ʌ�<�M�H�@^��am6��p��@w�p��L�����<�Sj}�G���@��oٛ�Ü���S����],
�D��%h�j4�%3$�Rb��f���8����H�?$���ww]$>��}��`Ὲ�������1�tdcJ�����y�+-w�˥o�'5�F鸩���������i�A�`~��D)bΉ�H�i�3�"B�M**m�����/-w���c������1�^���:���g;��Ns���lsؠ�iCTτЌ���Lí]@U��X��A��1��)�KԂ=�V�]21�H�A ����|B�@6�NJR�)�i�Q����J���6(<I��8�@��D(�}R�o�g�,�}�(��wٿ3���5���W?_����K�� ��/-��}�w��'�ti�}���0Y��]���N�ٯ_0�W��`�����=z�6܌đ�v���zǊ.��rVFJ��~��r�y�֒풽��Oy5zn�N��������u;��#@ImtKi�fzX�E+����L�*b�%ek��b�V^�p��<�2ET�w�Q�;.DK�F�2P'�Ϯ�jC��h?��7{ϐ��[����3��Sӑ�쯜��<w�Ұ!�j�LQ�쥠�"O+�3�j?��9(���~��e�G�f�U�m���]�='e�B�X 1������[�}4���W�ɞt~=�6�:.���bekjG��\�,
v� � �c���B���
�x��>��QZ����R	��T��"�'��s�=#('_֛,�A27eD����Ѭ��7ˌ/
��#3M����t�.B$u���W�u_\���p���_�S����������cL��3�iѭ "�e�b���>����V%�`�77ٲ"�@��G4�%��Y0�`P9��8��#�[2��uB��#�HR��)�ߺ�MsC��5^C��UYZ�INZzK�L�*0�� epHi�U%���\�[�F�*fFN-g��6h�V~�s볶F4A�OXb~��	Ո/��$�&|}5M��b���T1����y�ph�����xOu�OP�l	˜��i�����e�Z֢N˞��A��6���k:���]��)�|�5��$d��Ұ���H�&����{ǉ��.�E��%�.�B,z��5$��feGSx�?��/?��fn��͞�U(Ae]���i�H����p�tZbCJR���;��ޘ%B+&ȸ�<��p6�����Q`�WJ�^9{+�J��"y����X�P�����<�]��1��I���;K��I�c�OQĂ�$y�I���_J�0B�]8n��.Uޭ� pV� ���h���]b�0����|�:H��뛑2 �7�1/#@ٸ�4uq'�Z�k���nk�͹�#�Ôdv Z�D��s�kܔ���ҁ�BzK�DY�4:���c~}���� 2:�L�����H���D[}���,�"Dޢh�U��2-���M�M7��Nά�`L�ZxY��Y��^����uoC.�h�Ix��O��2ُ�)��~��%�ae,iU9����؍�}u{�?+��*��=)	�k��s�畎����Ӄ��+��\��XA����J���r#M{�y��,��H��9�����U3qC�F�CԾ:���U�^��@�0�B�@<�����iG��X�)O��0���u��a��.
�7��i\��S�f��m�3��i%��6�o�#畞��
Ef�{�Sc�Wm`�%ax��SY��z��
�F{���1!��Q�뾧ߐ�1�}b�?D�(���Ք�W�远2'��L�P��GTn�Е�C�Fh&e+�ߣ�&&�}��~|�*J �A*���M���/�"���x����3��� �nH��-���-S�R4�|��
���I�B@:]�?�ETe�M�颡�������flpvM�֩��������Ca=7/�����A�6�/Do�K^ގ�y�w�O�6��;׼X]�ٙvZ}�`b����K8�笶�E�@أz�=�4�wE����s�A�L�P��w�����.�=���W#1��9B�&�`^�
�?f2kD�s������B�[ ZY`SSg�
TӔ&HG�}�0����f��5���4O(ȟc�=�B1h�e0����^`j#�?�fB�j�"X�v1�F��
����+>/A�e\�J��c�*�֧�0�����\g�@.+��̡��<sw�4<hx�Q��ߧ:<}[5�.��]5U�$�0q�M��Y���
�G�H���;`f8����6�vI4}bR��bX)�4��"�.@��\w��I�Fk�.��yѠ���[B��оmA�a���:.�&f3�.�_�1��h�d�� ��j\-��?bd���8���d��RQ�/�eܖt&��ל �59��z+���5Q�1{C���1o�=Xp#1����ɜ��`>H����)	�l��"<��Tj.P��1;;|b&gH���B9�-�>k��z�<ݱ�]�d�>�������S���"�4y�!�����0��-�!U���y\��0��M��X��ʓ���$dd��]�q3�Zz�4l���fVR)⮻Ul��8L?�
��wF&�1���e{�$�T�YQ�_A ��Y3���B8|�I^:l<<Q6����v������$����zD�5�V�q{� �2�]�(���C+�*!�*����i�?�Ȥ����l�S��79�E�ɛ.V/�j1\o,~�o(|m�d0�K� �z$��u������P��j�Ǯ�X�d�; ^$���,V^� H���^���D��j�����N��"�CoWu�N�R/)�Y��s�`}TQ7��RM�VZ��P�7�g�:+�����t���-/�m�Mn#-��K�g��L�)����%Z�X�1��43��N�5r�lcx���ώ���S���,ܷpv-s
���yR�_�� �ol�S�M�������V�:nJ3t�'ș���P��>h�94��C9e���c���%�{��vOU�3#����h+��eD�ktӥH�����!���Sۛ�����3�m����T��?A�L��{��N�9�f�M�aZyt�u?�PAkW �n�R��w�=P.����&`S?�[�O��EH�
����Qs��R"O�d��b��KB�y�hh���\���~q$q��m4�Vl 2���y�P%�#yu=\F ���Ԏn� }��0M< ���� ]̹���ϳ'�&ٖ�w�iCD�O ��w2�e�J���ھ���RNj�U��br˕������r�`lV������vtW�v�83�`k���X�Ԁ��r�ޗ�I��Yp��)W����n���>-��Q���h�3�B(t���0��ftU9����O}kix��O�_�כ�A�×z�7a�x�����f������|��՞@l\j~������U&�q�S�ǥ^'�h@�b�*֦�Z$-;&�X�W��S��6�i�ٚ����n@ۡI�l�S��mޟ��2��qt	�,�LQ/e�nv�4���<g9��8s�Ud�O�S,$��Ν��p�<�
X�|;�D8t�����`�p�r�%��ﷳy/��v�a�yS)A�9/�]�����y�b�2d��{{dT�A+���3s��ˑ*�2��~2<��w 0P�-���;p�S��:/E��u�?]���E��y}τ�#���tp)R�_E�����ߖ�Na5�#֗)����������jؗ����Ĵ7^x�����$o�?&+�{�# ��Vރ�*�
�|�d�L!'f�xl(uEJ|���t�:�8lu~��s�	܅�;�ؔ؏.��l��b�gҜ��P\�� )�tDy����pu���|�L��+�QK}��4�E
wa���ap1	5�r3T�WNf�� ���us �7L��6�oT�	_G�6��\�Tt4�G���g,��Btg���j��B��|��ߤ��qr���������o�)e#�w��͐�&RZ��DB-�4!��]�a?g���t�AT�sg������Fq��%���`��K{8��*�G�*�vQ�7HW�>Њ@E8�L�;2�M?���F0Y�Z��.��|��+��ә|.�KVhI5�s�m�݀:���Ѡ��X�cI����rO���R��/mR���d�� V�jعO���R^��UWq��h*�^ݦKMk%�f�A����B��1�������8��!�3��8ls����N���a!�ǆnU�Q�C9�49l6�z�+�\8�����Xj,)�]jͧ�= �/�ȅF�N�/�Y��A^(���ʪW�����2ݲ�37���K[��fA��Ɂw��
��z"��s*G*���dK�b��]�)%���,���_Q��d�h�o��ݒ�����3�����4a����v�sqex���z��,Ր�%�7��X���z�Q�n���%h&���C�I�ժ
/q7P�Tc�a�5���R�0>��Ҁ��G��Ai�ۖD��.�.a1�� �ï�sS7�w��q�_���������W�7`�$�-v���͝$���4�͏�&
K���>ӁA>�H��*{ �q;�.�"Q����є��ҡ�]Ԃ�_l����y�F�WP��?4Z6������B:=y>��̅ٙ���P���IG���}��s�/�4$�"��Yma��l�r��=�Z���d��N��Ļ0��)�A�NY�sk�t�����>��&1����t����!�߻y��� ��u��F^]���T9C�)#��dLG�)�?"���a$d���ef�t�\���'b4ׯM� ��������#M%�1&��4�v�M�&ܫz0��;�l�~/b<��G��� LT)Lfh��o�O����y�#���� �� fj�%���1��B���*`��>3��x:$�:k���ս�;���7kL��#��X��
Z�j,Ӎk��M�H��g�e,�V������a�ʃ; ��Z��@�ۣK'���JW���� L�c�27�[1�U�#&I6Wz�^��z��}~�,7R����̿#�eE�o�w< c������E��A�m���3�M�z���^��`�\F�tJC�i �����]ӘJ} �J�a��1�j,'�q*6�P��FQkR�(j���EqY�~�X���ػAZ�^��#�RC��Ǟ�(����-�gbd��;��{,�q�^v�`J�=˱���V��/��Kv���'�H�~il�:ni��5���a���>���ǣ6�����T-�w�^O���y0��'߬�𣜌���]���Z���r��1��~�4��J(�\.Ĕ�#�xX�9�_Hh?H���_>�r��Ei�g���&SJp9[�F��DM���l�iN��`���Y[�^\��	���g�(3[�m����!g�����ȶ����&���I�*qD���Y����+OT�Q�u��F��"��v�v
��Vf�+��kL��P������	pp�,�s"���4��9��k۪<�#S������P n#�oϐ{=&�j��Zb3���1o����I�飁Tr lAB���K[5����^�lu��ɸ��u�>�u������r�H����������~�W�3���M�e䵊���[I�q��A��yb�#��gZϘ�K"=7�iž����ۨ(3��R�%�~ř�*g���F�
�РZ?���)�Z� ��o=j]�c/&�e�0 �>RQ��H]'�Ґ_�0�zhN�͙B�(a�������wQ�p��rN��[�=��9p)
�sP5�w�S6�.��<T�ӥ&�C���/Mc�d���#"�N��L��O���e)�7����1��UM��?-z�O���DϏ�ؤ,kx�r?���j�Z�q()��`�m�^�u�
&<�Q�/�� ^h�V��dS"���&��zk�.�l6��	��BFi�i3[Z��`a�t`�y��\4�✉��Y�_"�	�R��{ʹz�^���7>+�
B�O_�=	�I�k��?���
FY���C���@Ÿ�j3|�y�+����^:�XW����jۧ��0�@��s���|g�Ĉ���8�=Ќ��x��l���Q�,��2��i�%������ս��+�1K.�k�7G�G�M5��񔀙d2ά)��hA�/�e(�,�gt� o��]w��y��h0G?�{���m��*��m�G�Ɛ*:��9K|�7
����E3 1�R�|��c���B�����w�LPp�L���%�W�dR���	����P�E�#��L󵦡���d\�W�����EH���+Q�B��3dUO� Ұ�E�,j�O�*Y�z���v����T8�]��n�)$�v��Y;%�b����� Z�eC��"Dv��h�Z[
A-A]��������^�4�|�?�G��5����}�$?4md��4?�hy� m����m��<h� F<B7���4��g5�5չpE��D�׈�-�ׄ�9^P����l�ϚFQ�[�(�6�s���'SGj�T�C��uZL��>-rP��o.���ఔ"�>��=)|��PƵ����%f������(5(�h^�ʕ�S�e���{��������ў�L�ki��~�f��+
���<���E�b�;��VT����N/x8N����"jK	���:��5�3��i��K���"KyW>>��9e?��HZ�Ж�Io	�DڔH���a9��5�;�\C���z;/F	Fk.����ۚ%�޽Ԋ�@e���_�CHk��= ���С'y�S����l[^6�w�@g��`���֓�Ҥk~V��_��������Q��?͗�>°���4����Q���V����(F��	�fLA�u߃�R�U���}������bF}7m��B�s>K�_X"6�<V�a���9���fPA��eJ��J���a����D)M�� !��6��/Q!��3�C�u��T�y1���򗂙I%�c@���i9$4iFI��f���t'��M��B+a�c��.��I�j>�sLB�8�V�܀���y(�/�3,��2Hf��۰��d�8� �����T�d�e���H�����;̅�([6$�����u�l�v��f@(I���:�C���	�*�̮S圞���B}�ù���f9:7�t~�3	j��c)���v��_ll�`I����RdqGz���[<�z,��+�s.�G��n��Z3^->F�%H$��l���'�i	a�N��mڴ�y��o�4�S��벯�ұ�oT0�^N³k���!����i�g7Aw[[Xy��oͲ���^A�נ'{��;��I����I��a��Ŵ�k��b�g[T���BNd��8�c/P�j�Uc6n�,�?�z����O�|�J���35�8Lq�r`��������lbI�?�*E��6] 9X%2��kjwo
<�sƈ���t�����ܻJT�%�;\+���`��H*�ꪾ�|Dx��W8�6 F9�o�*1�I��d4�a�g��i[�����^��~.�?j�@+h�Y
��رD�ҥ)$I���ؔ���������HY󱕖ä͵�svw-��2b��#{y���vѰ.rK0"�P��6i'u���I����ߵ�KD�6Q/�'�����լ	��
��H�����
]{�8�K�
5
h�����3�|N�
3.��ՅA�n��J�!�Y=,�LbTp�<�m]?��nU��)���Ҫ�F�Ʋr8�8���q���
SC涢!��RǤ�M�K�B2�S�.�(����ڼ�-B������"|�u6H�缣��cT���z����5�>�7Me��.��\�������H�u2��U"Ltb�
atID'c @�.^�~�4�����s�&��?�#A�]��O�l��ʹ��mr�vt*��kc�����OB-s��4]��J-���ʓ��� ��@ŝ�}&��x�M� ���2(�ݏ	pǪ���0y�]M��)a��)��(�d��4������ۣ��.L�GQ�M���9	�7�"���H��N�bN�M�X���^�Z]�rܐ��nݞ"��u�%Sl��C˘�0+&D|$D�Ì=����*7c�"=�{�GQ,>'R3P�f�C�
ΰ������j&��iۗm���9!�Oɕ�d{E0�cR�[l裕�x�>!�<��BB`N˭�����,p��_?	%�iOL�tJ����ōD�%����:Xΐ�l�����W�A�KѲy&֣���Z4U^�e�߀G��e"���h��0���>�uy͆�������=���_� �\P�O!2����!�$��B].��-��Mv(	 S���g��Rv"{\[c֯����s�&	շ����=��������+�<�^���⿈m4	@�
�#��o�l������,[�$V� .+���n%��lcJh�' ��Rܨ�n2�~q}e+��f�svA�l�L@ʃ��B�?m�4��`�c����Ma"���ֲ�6ߧ�>��{�D�)�7`�=�I}өd� &����}U�3A�N�~1/�sZiDH �K��̽�d��|�}A��J	�����忺�z���UB�>5��R�=�N���l�=��b]����CL��CZ3͒\
c��|u��J64�H�px���4���Ζ&�B� �~�/�DN���Rhv��U/^���(ë�%�WR�޷�b6yg�����
�f�XA���j��4@{W�3;�9#�YfS��2m��t|�;����
)&��V�0�������K�9DW7���p��<[���"	��{���~O�t������{Z�b���z!Fsx��y3�D�D�L�p�U��ޗX#jG�R	����A��Rޑ{�)� 7���kk�t1��� zƉ�����[��w°m��H8��M���zJ|�Y��޶��OjgXk2<g��kdd� ��S�E�a�c@Wc�9�>?6����ݿ�B��D@�m���;�֎-��m� �qLš:�l�O߰�P�[�����]=�XA�x	Ru�j��̲Ez�?�CI�����b�^9+�fJ�g��8PPJ��Wn(G%7��쏠V����Q�э�(mZ%�('w����>�Q�Nm]5y}n��������ǥ���l�������a\#�ՑM&��dPXg��Ro�1Y���?��Ď�甤I�|�{�y�>4p��R�T]6�Sx�S���|��1�u�,��h�i�P�8{��$�����~mf�V�~�
�@�H��v�������m������e[
����Ak�}tj!9W=OK̆�Vbyw�}w���է�7=%��i���z��x�bﳖ�"ƕ�6��|����,0]{��w}h��9�m�oh��щ�LpkS�'CD���"LS�����|����d��3��.L�&��_��8	vL�����%�Z	!��l�n��i�k��M�UEGH�I<`\�{䥤��A�Ï.����F��C�|:�T祂ԡ)��&��1�࿹Il[��cG�&��?��8Gky�����,U�^R"^ȼ��&����r>�إ�,uT������:�i���1�d��I���=ĄWM�L���2I��P|�n�p���O��Vޘ�|�O�K�O�V4��4׉�G@���$�j�ݟ�z�!@%d�B	�*t��.!B�p0`��}�'�kV���m�ø�
�
�܅����,5�A�7F@��j�EQ29� %"��M��g0�g�A<�H����/`��/Cq����r"nx�cI9��4���l�0nrKQ�j;��5m��a j\��& dr���D� ��_l���/���Z�v�Ɓ��qxulr!@#k�(h���򥴛�Wn`�����[�/��&�O�+ը��򡆉�h�_��l��u?FH�#�؀��:�*��G��G�ǁ0`��H�I��Q� ��+G�@̿�h$�E�Ȟ'X�f�A��[��2��g�IT O7=TP�z�e�C,��P��cr�r�F8�VMˁ^���F�)��+6��1���+�z�'��Ӎ�D�7�X,n@��o٪�u�D@�ޡ��U�_�� Aa9~el~���v��noI#0댢1+�uس3�+���n���k#�O�������
9�U�?HDaw,�K�
_��/Rg�M.=�*��/k�s�X�Ke �Y#�X|�����Du2��"pfO��3L!���@7�J&�P�Gˆ���,�︞h��۔�[Ƣj�����h� �<�ܯN'4�t�E$�a�;xf����G ���9s!$8�ט�M��E�I<(t�U��mEۗ���qKf^�� � x����G�1�"Ԇ�����Y� �'�{4��~��*fx���`�g�5q���:�RTpBG�����K`x8]°d���{�'���!�S �s|C���J��'�9N��cWS�l�O�Ys8��?o v�();�l�.����K[��5C���QK����gS�L�����$�C�vg���S�#�(��o䗷"��[�����Q��&�{,�Ջ�0*D�E	��^A�@���as�'��+HPeI7���ȨnJX�lZ�Z|�JY��T��{�a�6�(�M� � �#˾��Kj��@'�������!E����^8I?���xE�����1-��;�"s�<>ٚ�2m��� l�BӾU���Z�O�'��G0��j����]@�z�䴦I�κ3��Ȣ�n������r_^�7S��F�@���!��A����\���M�O��6�1��?l�=s'�e�!S�#G �\VP�&BG{vշ�Mn͝7�ś�+�
N"�ݎ����W��(S�B�{l�`�w����uK#HðJŔ�n�1X��m�5~4y�\G/��Z>wS�
��.�O���	��rm��Gꦨb�`R��f_��x��]rs�e�����K�XJ�R�j�;tK�O緲Ni���>�i��U�8�cʕ>��Kh���e��RL]M5Qm1F�DB
9�`R`s��w�Ù�n-�����x�;v�s��0��ЯX_$S*ڔ��D$��}����o9"��x1������Y�1mPu����h�ue=!d>��JR��pN���*�9����5i�]E�ڨ�����̇�\����J�Sڃ6�����24bEڔ�R����a?����gi�f��_�����I���E��=b�y��r50Ms�������	�N��/rXrw�'H�W"�Z4CK�O�d�^�����Y����1�(�>y�Q��B��$@��S=�x��2O<�̙�	�L��O��3o����״�w�1�N��DMok�
�W��Q0�T��&d�o�,��{M��R�d�=�����~?��{��0q@pg���h,�|�z�0�(p@*�l�;��T��-����)���!�ԫ��
ޏ�=��;#��UꞰ�[�Q�*+C��ԏ�r��'��7?[,�����=8�p���V�����%B�ۋ�����`��ì>����'�"-���/4��`�A��*	�G]iU��e
)v�8ܤ��io��L���amR+�{R�z�D�;@E�O�X���qJ�R����1���@��L�0L�-�'ୡx	h=l�]T/��
,���xS*�zb�O�E��8�����l��3�4����͗;uV�A����m/=c(q��X�.��U��U��;`m�}�]�: ԕ�i�O`�f�y6�03��7jo��/�G<f �_����Ay�۟�_�)��I�qǩ��*8�������FH�ߠ@�'�Yy_ϵ-�g�d�)���a MCY�Ǽ�t
�_�?��i	 ~Y���{�Ok�"dVLq%��e���-���û!$"�J�%/XG򤭚J���k��'Fy����'�f?��!�L;�=L./���N/4�[�����&-��?utb��W3-؇i��7Ď	ǉ����Dx3�ʯ��kI���޵��)IB�墱Ļ#�c��->a͠D��ǎA~ڞ5;r�MH��b�o~^�͑iK��E%S��C��U���5������G��B���
	��sԁ�F�|�/�I~�۫��F¼��H�ܥ�ۓSg$�����܈�uK���`�ة�>�i�l�����K�UR3�@�*�`��7f��ֱ�^�w#� ư>�K0�M��d�����$6�y)c]�W0���?c�s�ȐF����}Jm���n����>�E.T�T�lk��x��|���hQ8Dm��O+zٻG��q�m�����,����
����w:lT���J�݋��)+��9vɍӯ�v�Yzzu��q0��ͱ�n���bx ;�=ֈ�Ao��b�I�ޘ�1�V�����`���պ5�����혤z&W��ʵ�T}��@1����C� ����2�,G�+2M������7� �zxs�d�1�:�#^��`�����:C��RS�:��<���f��6�=��H�/�x!L����$TD{xӕ���IC9f)�h�u��`Lq���p'��G4�4h���.2�8�jTx��\	�=_]���**Pj�g�� ��h�88ޭ�����8�L�{����������R�b��#�4���Sͱ]��k�-0g�n����`���y:�õ��m��y=��Ӹc��P;D�x�=���B1�6E}�W�]:D��?��!����*�L�H }��#��v����A̦��tp%��]Gd!=�<re��@�[�Ua$ ��}�η�r�y�d=l��N���ԼS}Q����L�lPZa��	u3S$�l�5��SGP�/˫�=[�NI��~-B����"��A"&�}ռ�WN,��#CB˚9t���ß?t���Z���iI�監ߏ��K�d���.h���{=��3�3f�^�d��0����m/X��:Gl&�КOqY�A%ҁ��e��`�"i�]@v��q!��+J��g8� ���� 9K 6���Դ�N#����g���ME&	��u'*vx��0�����xK*>Ǵ|�u|P�b2��l�˺R0AɡGj�$U��p�[I����H	5�v����y�u�b�'�1u}�x���nzL�'7�6����C�fF�� 5׻�G�H����<φ�]bf��P4��f��:�F�H	0�;�;��S��3��A�RK)��6ߏ����p�� KK1�&���ޅ��Ed�����v��yH�Sx�5�������΀S|9�=�kY��rT����o�N���Xi'T�Z����1%��
+�q�v�LI`���Db��"��!<7Z`��(�k#�������6�7�λH�*%�z���?a@���V�k��T˺O����^b(_�jڠ�����T� �`Í�`ҝ-8U� �(�>��B��~u�%����*޳>��y�#qr��J
��c�t�u��
����帍���@�z�ʝ�p���ND��:��ܺ���j���J?��������e'[�n*��]0"j���!�s�s�J�m+�ؼ�%	p��Q�Yz�� (����rF)F^O�� ��@"ub�r�(�!��tb�U��������� El1p��z����r������v�J����A���������Fёk_�|���	a3S���	At�"�Tl���>�z�/N �V�$-.Vk�u��	Y�մ��65��ƍS�q"�}O�I�l#�����mV�$���D_`	���3~�Kf��Z!-w�K�Ed�㈡F�=��ˍ.h�X;�$�ձF"��� �!5�ߗGSPʃ}%u0�]�T�W};� R�:Kp&ps6�-��.��a���B�sbI��;�e_y�V$�M�mA(�Y�r���3oc��b����o=x��ܮ͍\�����i��CD1z�h �.���Z����t�}mc��2N�unI�:�	�op����TF��|������I:2��B+����S�\�S�V�`?]AK�_���ϯA/�1�U׭����$��_g�gqZ!�I�#�;�-�T��Z$	]��|�9�H�t�I�H+�� ���r�1�E�^lgٽL'�w:��b�<pG���I��m�؁�d[��M��/�z�=�� ���o�a>��6���X�����d��c͑�xhg���W�
����?[M콜��u��E&� t�p���"5<)��:�=�Fz0��a��sn&�!��]]eFQ|8�ua��Iz�շ���:]]�N<�ѝ%Y;�L���PwIuUX�]dA���p�����2H��-e�F��*l�q�)����(��3�W�zt��������RC+ut�C�*U�jZ��;Ytv;���!2�E7�C��جr���Z�ݾXl���￠?Cl�%v�����h�v�y�/�7o�"���q�H�P�.��F�-��hP��C���#H�b\u�Gr'�բ��\`_��� ��Ϻ9�Q�z��Q� 9-�`�����II��H䁑h�Y��Mw6q�F�<��z���ǪG����m9}T��<C�^J�CX����s��o�2` v��:||���h��uZE\�(Ė�W���f�٩���wD�n���gKU��4C<���=�x��jԟ��UW�jk����~��$4�T�P�Ddc9���K�oո�آ��W�D�t]��~e$��_�,�Z u9M��I!��pB9k����b�B^�g�E���[F��O�sXT�gɌr���"5T= ٪Y���&�U�3
{���lF�6�U��+g(����Vz�m�h�6>+���XK%�?xg�m����>s�lO���^M�0��ހ�ͽlmp��Ol�<��tw	r�A9j�AMm�]���n栉DzK�R�ְ1�VV��gҙdګJ,Ԧ­jT�JP�M�K�[�(��ם�4Y;�fGwwN[U�[��Ri"�,�x�|Ƌߓ�6��D��U��ŏZ�x�p�������*,Us��L},����{�@ܦrX�"F�r�q��ՠ��};5k��ٓ����mAzH�85����p��%���`��Ӡ�U�B���XQ��ˉGn��JJ��`l���x1y���Й��s~�\���w��W�bH���J�!��1 ����ӈ�je�0�[�G}��:�����G �
�e���֘�Ul�~T��
Z=Y��f4q�ן�݄��,pDPsߝ�����/{�.t,��z��*HqB�c�z`� ���J&g���ԧ�-�0�FP9@�^.�xn� gV�>F*6���*��9=-���]�����Bc��q<��
s�1����;E&����F@pTٴ�೾�ј`:s�
��7��^&���[� ��+����/;�dS��3K����9�$Ԕ��A�C���Ruq?#x���F����Hy��(��*o�n^ޫ���O�����d~u�-��Kޟ�i���S&OZ�a�T�����gA��>�qC���.*H�|3]vkt��F��j�nѽq�ͧ�-]tb<��qi&���t����	D{�	/Țݒ7n]�^CF+�<GQ^����EA��.����m$�pU��I�
��~�],�}`�A����A0-�(:���8�o}�I��8��ǞO���$���l.Ws�ˤRQ@�RV[��ո�"=����Y�N���F�lѤ=hoD�U�+H����\s�/��a�^w�fԺ���Kv�<���쉷?v e�5�^?��y����A��#r��,,(�n�ǖ9ԒS��I�F�N^�b*���^��Z\���0С]��D����2��A�*|�dP �S&*�f�&�0��H���!k{}� w�߂Ti{��5�\b(���ct�ꐐ
�^\�=��Xq�(��ȅ���,cH~&��X�����C�R���<��o���v "kw�W�*�Ғ���VF������j?~:�h\��?3e���$�)�lH���~�9��
&����[{�^�i?0uu,��tU1q��3��O��}��4�գE�GJۑ<̺�b�)#�����S�\���PD���<���ӶY���� ��#Gl��.u��Û��l �)���@���	��;G��_�kW&��{�O�Q����nf9"���>M�VOnhv��w7��n����/q�Yֺ��8���4;���1(ԟ�f��~�?<�Q�=��XԒ	���+v@�P,s�`J������Yn�S?����(��&D8A�>��Ff�(���1A
C/�ߛu�JÆ��a'XhM��I܀�ٰ8�O�,-a����;}�H�U�\��YP�]4�Bx�ʛ񎺛�����r���y�w���Z���^�x�͘�/[V>��@�$�t��[RNôY�[���F�xP[P����?X9�J�O�W	���M(N=������	Z�����F�+��e�u/���'V3�U�d�M �!mq���eT)�(,f�?��c�lg+�4S�~I<��p4D����A�f�m���(�m��X��ԥ�/6$��0P��JE	��������p���Vq����i�BNy��G$����#�zҶ�s8�Z�����^���3g;��:�����������ֈ%W�]�7��ZZ3�*\B�؟R�]��J���R�Yj'���A3��%<�h�ƃ�s��R�j9wv椌|YP�{6'��M������	3ÉY��reւ'��!� i9a-�Le�~���b��,�Tk��J$@��-���/AC��bE���>��YG���s!|z��u�ٞ1�1��n��� ή:܅⻧���X��+`�7�Avll)�Rv]�J�̐�ɩ���A �ݏ^q?�p�%+Dp��|N��a�隇γ'վ�.$��l�j�+�����*r�����rA��֙��í��X��R{A��±Ш|���O���EpopW��4M<�h&�)H�0V��mm����� W�3G�=�P���`jD�/f���!>e����IR�dH�`������/�X�Ƙ�&�{tWȭ� ��4��L�؏�����cť��n��uO㐔KP���r.�H�+�G4�)� �i����zKjEG�{��X<������7L�_36��̔B�w����k>����q�~�A��L�g�0�ւ��+N�/�����P���bH�K��-zn�Z(`�_�-ʶP����4S��7Ȝ0N]�q^j/9W��E�5�C���k�~0r�����rD�z��OV�k�K�%�l�5!ّ>RL�fuM�w�����]�dѻ�XhB����	���Oh��Ů<=S�ݱ05y�O_�y�
3�*��O�&���J��5�:?�'��_9�H�-Փw��#0��@��G�����CMM� x���$q���
�}ƥ҅�)���D%�Nͣ�i����<�V���ݑ�!`�~&��,:�`�3?H�E&Dm�<���rFН޷辕��k �����.y�3(C���T�''T0�kuJȅ������ط���/L^�R��n��{�Go䔼�G"��/zc�=xʉ\J<�A���j���;���)c́�0`�X��Jk�_�BLW����ybm��-Hn���\��4A���Po<���Ғ�G__.@����)Ό�����@�m��h��e@�+S(�z����3�P5LJg��.�K��s�T����B�G%�vnmC���a(��?�ل����!A�nN��{��L������0A?R�˜�?!����X�_�4ΰ�V]w�c`y�����`>T8͐�Bmֽ?|����K�E`}��Jk�Q�]�|�ul��YHc��h��~�毱	f�$��[Ŵ�Qt�ʇ�������!�m�!I��5C9{�
�6�'<ފ{*�+���>��j9l\0�jf�5렏_�I�M`�1\-���������vva��ǈ��r˒{1�I����c7��S���Fj~�MXs�/�訮���Yv�cm�M��:(0�c��5�5�BA���y�X��A�<��u@~�(��\��������0d�,��[u��|��!�<P�Rj�S��\�E���gLv�1�m����t�~MVY��O��8E�zɸy��@�2Do(���̽0���rhP-���I)�{��~�c�x{�<n���sN �Q����郪�&UR)�_Ɯ��/Á����v��Kd>�/H�
i���ȩk��/G#zm�)���������u�,g}�L"�.�~����{�zf���Ȓ��� ���N�3�{7���(d-ɔ<������,���)�]&����1�0�+n�'�B��䑐>?Ua���HQm�B�k{D�. \S�����m��Ʀ,ͭ4?�,g�Q~�x9���M�Q�XN�q��O�1���X �L�2��z����Ui��d牿6���{-���&>��z��Eѧ�����޿OQ>��l�h��K�K�h����Y��O���Ԣ��FTcʉ�K��.[�����Gj"�G� ���Ig���]"8Гc�i��k,qX>![!�xM�>��X�+��	��!B��̯�M3����E����T�X] '���DQ%�>���"&f��LI�	r�kď�zS��凞���˗�uDHS�4��F6�"�U@�L.N��|�oJ��M,9y�o_�5�b	}�qN��nD�Un���:ް�h�+�Ib,&C�r)�Z����	�f&
����_[n�(!��!��D��'LAF��8��P�0	�޷���ѝV\S��O3 �)��)^�Q��X��7[���^�Z ����5ǩK�&����y>E���1��Yz��T�'�%fY��w���qS�J��0��Ɨw���&`�N�E�S����Dk4���&��U�]�� ���v���rD�Ĝ�1�5�Ͳ�X�cuB/�/�����ķj�V�Ģ|�,��ӎ�I��ׁ:-7�fs�N�%�YaԹV��B�RU�ɾ/>w:��J��<9W�d�ҘB�=�r�=��`M�(�*��1����~'��_�aG]Y�ZH�������Yi��<D��iw���W�&��'�-U�-��t�3���n�V�Eض�q!lC�<T1p��\�*��p�⃪�^qE>6������-�6Gx�����������/�t�T���FaR`��/��Q��W�l��O%D�tϢ-+�ɪ�mؕ|�A 6Q�^1�ͨ�!(a ��#��Fia��Z��:%a��gC�Y�����-�KL��p�0���}%��hnX�d^���5������^@�2�]?|;��Avx����ٷ�]	�Lm�}-}��(�4Ox�k/j�I,ه�L��_��3�`�|�g�[�wT�狆-;���^�U)��4�8�]��EcԆd���1W����-�����L��l/�!#@���Y}m����x���<�r�~s���2~ۊ��x�/vo�+�JT���gM�y��3Й��^SrДLӕ��B�21S��m�x�E�:���LF*<J�
�J��,;#}W����xVli³���Ŏ0�^�:���7�9`�jL�>8��#��9��B��7����p!˺�-I�+X/�8;�B����^=|H�N�����R��R9N���-k�
�.�� 'Gd�r�on+WVHuH
���x����Eyh�sfO�Jc��,i$2s�X��Ǽ����&��Lu흕m.#�o�½'�%�h��;1�0Ce���4�MJ�ڨ5�і��k,֊����̭H=T�!�_�N;z��{��� �z�`�i�	R���"n��z'˲	m5�[CI�ʡ�?��g�s_A9�%ݰ�򪁞xI�[P�^��6���~֩ɱ��^zy��'�
e�p��2F��XutP� ���>��äC��@���Qk��!e[x���c���J�ܩY��H���ͥ7���'�`R�~����,f�d ˺}���&�sa��1�!/5�G��៪����7�])%_!;��B��N'��:�D�mN�'��3g&|��@�(�<2:��xN��������~4��p9UU���I06G�KRUN0�:��k�]�B�$˺H���)�7�R��L��UPei�^bq�
��@���0��o�$*�yӦ3����uF��K`'��Z�1��Dh�z�Z��䴶�Z�y3�RZ��*u�gQ$£�b�n�����\���Q���jѰ�C""<Ue�ѵ���>��7�j��׆5���^���zM�2vD���KK�4o	a����~��a�:���'�p�ej�͂��Gy�݀��PRB��AsB#,�>T1���:{/cQ�Zb���­y��O����BA|�~Y�Q�\�x{;��A�]�"�`���)"�+� ���,I��%��*�i�y:��J���-7Eʇ3�R��]l��~/��}>a
	���@'� 6>���o��Z�������2�?��>�썜g[,E�!;	g����+��2����%Z�|�odӹ���sg,�b"bO����5���ee�R+$~�ݽ���GGG�>_D�]��PEb�1/b6�S������I۪(�_�����3L��X�.C	�7�=�3��-NXCOl5Ӣ�ۨ���ЫW�.^�cG�އ.n�=���łu�hP�}�H�8QO���_������n�C:�RYrÚhA�A�*��̮l��;T��vܡ˹�fYznՅ�o�8�T�N�v�"3��&9�Z������]�x2G;R�<�Q!Wr�9!�Ry����b^Yl�������Gy�tH�&Mj���u��g7��R�6_�h��2P���*�Q�	q\a�7�&g�9��*�o'���%5@��#v����~m�V$@����b|Ug�����՛k�6%�j�[U��M�iSv��?6I{h_/���2@L���5{��y��e�	�o��NTC��D��2K��N�ؾ���knL}{�\���~�����Xk�b����s��ݭ��Hc(E���I��TJ������m�غ=1JϿ��0R�T2@��?���V  ��X�*.b
�G~y��_�@8�z�B6��	�!א��oB��|@�?-�6�����%����z~W���(T��A�&a#���X�F�]L�0A<ra�$���!���1�ۡ�ܔ/��&V��Ǽ�ǵ�6�2���	�r��.�7�����mi����A�z���r��P?I�.'T���������}��u��ϞN~SI��4��MJ��hC�ȯ�g*��w���V��Fm��ug~9�(�.�a�o%��ԡS�������!��%D;	��{�A�r��'���� r<��� 
`+�#$���Ѹ}�&���@Q[`��0�Q�5Plh�_"ת�u�
h� x7��ȱD�Rh̀�pIB蹾�4��ͻ锲��楝����X�='NP��t���;S��������n��-I���g�>��߾w�a3�l
'N�cq�V�}>v��[,4�����4P�Q��
��*x�1�r�T����a.��fNu&��;��g�Л�Wmg&�F�����A��Pqt0��6�X�yπ9�$Zo��u��6�,B�-�ȡ�����T���.2��yh�@���i�/ �r��;D������a�g�I�@`�k�9)��Y>]ZaXLF�$�������n,��0�^6�W��9�d��IT����4�L;Q��,��{��H&m|�bِ��tBtp�[�c�J���sԊ"�֩\]�w��NW�.GQ�!:"�t�A���"6��ԡ`}����#�)��
.�D�ג�[u]w�.a�!���e�>x�Pf=/��C#\�����fr&!��_q����q��&%��}�	@�������f�E�/�'�NlC*���[{S�Qq��1*�=�E�w��x1���E�d���3 wޓ�/�]��S:lU�Gi�a��cJ�_�@�J��+8B |��?�:�d������Ӯ�A��Td��Ga�	7k1)��$z���aK	`'��k��}���<��'$>���%�K�X�x���>Jxo�+"�S�~�ͧ{U>��5*%���e����P�f�jH�z�|�0^��d��&�����5�)�����S�v*��P�Kx﹯��Vw*�mK1��"�:�2�K>�Fb�yE�1G�F�\Qb���� �z҇��L*�J�n��� ����]����W���P����-��ccO슯(�q��f6D~��߬"�i�ɂ�?�~���)}��
�F�o��z2�?�I>}��/�l���D��WU��h�i�2��L�������y�j�Ks����g�u�V�U�A�m�v]�꧲rt��^���	���j�K��
S>\�D����#W���R�iY�kO7��+R���[!#�0�t�p�M�����:���xHǸ16��u�o&�$�L�dxL�S`_9s�+��^�$,c���z�/6�:3�)���쾖�56B-,���äF��e$�6B�� ������K�LU��z��'��aG���r!��������h��p�)r��y�dl�*l���k2��������_��Ux�-�2L�4y���+�����7B�2B��o�% |�鄼�4B�ǩ�\C���ô�Wg梪\�D�g���Wd��J��̎�p���><��Ba�ź���l?�ܙQ�W��3m�v?>�*�!Ο�@��*?UÖqYӎEABG0}<�~��:���B��?o #��٧��3�D����$Mun�*V.�Mv�$�o`tY���5�Y�0b���n�M5�d��sB��醍�M�b��\k�Ɂ R-{�*��m	5�ӭ];�=Ԛ����~!�-�I��J����d�!�0�B�YP7��y}��)�D�#��`嗱�i�*	���,�qG���S!d��U�"�(/�at�KX]D%U��l��-%��mS�*�O����ڱ��q�p�|?L����#�gQ$w�ZV�N��m��z�{g����:�3��y�]��\[&���C?���Z��<��Xj��0��)��biRa����N�2����Y�z��,��N�Ոrm~2d�h��I[‚n$m6�ʳ�O��$�lW���;�[��h���>5����>>N{��('�T�� x�ĸ���ȁV�����1����Io;","#ɡ�h1r�{I�2��b=
��W���lw��u��|�K�#�qr1I�h7�@�)�״�F�# �B�D�8������l�l��,�[���.&���d�ƃ�ퟓ�d��綖��s��@��&���Ӑ��,�{���<`+���y����B�`�qj[Szu���p='?����1
�n՘+[d2���Dt����}��W�����l��c�'�N�m����I��ְwϫ5��3��TkM�ʅ��X��#�~�!+o��Z"��[�ߦ�8H�y5&�{�d=�֗a�(��!��:V���X��y59|��@w]vK2�q3�r~F3�9��{�&��LW�3�����lf�T<��?�D�y��(�\�p���L>����UQ�sw�}1v7��ҳ��B�tF��<�6&K��y^(4U.q�p��:�㠊zg�,�H�ףL�:�.X���O1cR|0:�<����Ұ���E�#�l��I���s[�\�c�Y��� K�A����;��� a6.ϵQ9���~�p���ﻭ*Q�rmԅ��
�mdC/6[f �W
rg��*պR�k��5�6N����I���&��-S��>q��0���a�JN6
�"�����2��YS��،,K��!�A���'3,�,㒸g��Q��[�*I��+�Sw�ot��0Q��*��}�FC<��vz\�$00������Z3ռJR�&��-�B������C�X䎘��A��x~�S�2K����I��!�B2﯊z�	f+�3*���j���LH3�T�s�f���H@�$ϐ�����"k��^"����!��)��`#nU�ؽ1����b�W��J����-%�2T$�(2�u���Q;2d�I�!�N�TE���Pm���1>K�����?P�U��\w��d�F"	d��3#��r�s��F���A��8����
�p�v-� �&d�m@5л���a�~eW��n�Dx� � �B>:����.CAp� �h�ܶZ,>�I�- �5ft��	U��ӂl���FP�0U�C��VX�/<G#V g��|�m�~�%s �[�y����S:"���Y���?���Z!r���Dq�Ke����D�ذ$g�,�{*:q�9���-;L�(i5Ps�p;6�_l�����~m?)�fo)Ѝ�ɊI�P���2&_ح�uzX�|������oC������G�?�'�fb�9��tǵ�P���g�
�W�|��6�(}V��/��5��4��If��7���oV��f�p0@ �S�(����Nƌ�I��o��dP0��=���垥6a���h��&�ID�gP�K �u�yc�#���¾�����`pDo�.(0�H7ڙ�X03��Q�����H�K�F�Dc�E��k�/�ck��x���쎼r�!l#^c��+��!>���2�=/u��;O
pc�q��U�4�G���&=F`��ϭ�T9�@֧��,�%wAg: hE>��'�R%�6�U�5����r˲m�����iv�_j0/(FQA�,W�5Dz����_),���b�͙uy�=�k���S���� �(���鲌g��Z�+��4�m��T��G\K��_�x
K}qL�d��|����\wRU���7[�T�Lbq�vF�a�0�u:��m����BȅJ��'	Sw���K���������B�&v���D.X��4����޼?aI4C�M���D��"��s��%G���� �B�x_���;�N}����%���e�rmC2$����O��M���\-�6Y��6�GVEQu!�M�]��$�s�%���d��7�/zpy����K���ލ`����3����Юo�}�x�:����8���c�}���5]�$i�#���f��\q����H^\)��KG-ao?V�����f��;G��3����E%<��e�S^�0�S�٠�5�F���Nɮ�qZ2HE���4u^ʛ���(���s����B�4uA˥�0�?%�\�0�;<L�Ǖ|ő@C��*(כhd���ޡ�ᤙPf�]�1�맰 �w��"3�
������ �$?4�må6- ?�w��(�)P���z��q��Aw`�0��kA����.V���_ ��>A�[V����e���t���i�G�F0S����W� �u�� .��&�M`� �4�S�Ia�G��C���y����q'Ol1��� }�@U����Ct� � ��n����"(3l����D$IC�RB�l��Fc�I2�OJA�I�~�F3UQ	����	Z0���1	�^���. �o�콍٧���i�}����cE�^�K�p�����J�V�\�E�����ƠV�}��:	��'f����F�>�����$A�j�zzc��;�5}n^��W���z�|{^s���y����D��_#�� ��;Ͼ��j<ʪ��+:�N�G��u�K��c�'7���`xgc��3�������;JWd(!�䑅سZΗ�.�	���e�í�;���q	�	ч%u�-a)?�sρ�v�s�����ۀ���Iv���!6�+Ls�na�[�q���v��O�I������ �����0$hm�9�{B�=)�7��Nc�*��껿�u`���z�9�C�N=M*6������vsL���R@�iGZ�M�F��#�d�ҷ;��ε|���#���"��ۘ\�u�����f�&�b-���m�N4߅��(;�[݈�� ��.��P�,,�_���� ���O�N��3112-�!���i��9ca��>�h�1(f�uQQ�v�ڴ��W�����-I�V��H��J�QP�Y'.�8��k�����i�#���8!�c��^P��'oaS|����3�ŇF��%�V�-�����l9��}RaӋ��R�A݆�����y3#�}�K��4L_�ܝY5?��v����2�{�$� ��P
��ȕ��͝"3��nј����V����y�����gUU�"�9��&db�R��P�*i�4��/��(,�U�d�%��Ě�*P9�QQ�����Ug���ٳs��+�_���r6r�C���ňY��6�^�v|>����x~X�aը0���-Eq�a��Ƅ�)�'���ݵ�\��Nhr���ַ�7Ԝ�G�>?a�e*G�S�j�����;��qq-�
(Y��dώ��D�s����Y8A-��������G"'�.l(-]jϜ�2�q/�됰�o����4dԑVvtB�ZL9�L��H6>8���Z��͑u6�_�l�DC��I���B2��N�[�-���kQ�p�7�nQ��K"����,��/�R��5��J� x,ݤ��ed�����kٴ�՜ֶ#�:$�d��|!4su@J�1W+�*uG�E�P��HUns湽8�ۑAX�
B�����@ڱ����ZډO���϶�a3�]Sa���ks]5r�&#�-h�N��	obqC#)䥿�50f.����an
dx�X+^;��ZO�7U�8�kգ�!�Y�tCz�1
�����ׅ�� �$s��?#Q7н���)g�6����IS����2��cS�1C�`Z��#
@wM]�Y��xxgE�������vó?��{`�7؆h��t(�P�w�6�V�g��C&.ĲM��������V$����_D�>SL��"�GJf+���yM�)��`7��N���$w�t�c�����#G�"&�S7-��C>�O}qgi-�RƟ����ϸ*Q�T&H�kdӍ@zPI܌&�N��/n�;�-*��H��z��h;$�?؊�rL[/z��Ч�x<���Ƭ�v	x�_�]����!$�2Z���&kj��ho�V�0��qK���=�n��~�g����ÛN���J��kճ�ܴR��uT���}�_�$-���,~��?�_�����6sڦ�17�Ih�8������k!Ob	y��*hv��U�v�rh�C�<����l�F^�lMA
��F�Q�����20���T6y�Z�aO�7��6��L��q�V(�O9(3����x�<s��\��Ӄ9h4��@W�ѨU iO�j�z�*n[-��Ƹ�(���bJq�'$�>(��X8�'3�Fޗ�%�"Ӎ/^x�+�pKE�[kS���ݏ/��M����98�E��UҞ�c�j/��)N��ԚvM��ڈѨ��&�H"��&�e�b��VB͵���~fwJU%|���ר; �l����"M0�YT����Șa�����N�e
����Y�-���K�j�ayyV	��q���%Q���Sd_끃H�5��(��I����bF�)�_~�	����dE��I��*>eY�.2R�I)*vE��~�K��i{V, �Ǯ_�}y�?���������N����j����F�`�K,��|{P}�fԜ���8.&�k [�R�nϖ'�.vW�j��_�#^�]pbnv�(��WekE�������*�-�_�S��KeprS��zB�jR'���Q<����~+���Q'� �;��X���y
�M�nh�2��C���R֑��II�*��+T�1T��rW)�c߆�ڹ�(c�7��d~�G�<+�J����M]F��0��e}_��#P5~̪��V6����'�0�.�������LO�9ɼ�T,�z�/`�rQ���om�ph�5dT�fd���·F����Ň;���=�h(��@��51e���2�wH ����niy�3�����jƪ	����u�2�9.�*�QK(��6��n6i��25;,��-S_9�8y�q����/  ��Ɉ�tx�I�đE._�pZZ@�*g�>�
3��R����$�����E����W�p�^��~%��ʺ&X.��� �H~_L�ۈ܄��HD�f&?�̓��*0TOɷ�yq�) ��)D�3�.�?�`I��M�e���;��n�4�*Q���ͳڙ��"�c���ٲ�'���i�� ���,��E-�;ׯ�Ra��/R��5���Z�u�h��&�^�QVE�8����5^6�Th͡�M�t��J��J�؀yg8Q���FR\q����л�5�s��[�!�v���x�����&f��}DEy�<�S���?��a&�g�t5hYL�:����	>�.�5���[�>90hÑT�c-f�s|A��O��Yp�L�7\� ���M� ?�ڗ�%�G@��q
m�ؤ�,��6P��Fwݐ�~?�gϱ}z6����>��&���$��P�H��#+�]����B�2A�:�G�!�j�y��a1kv�V��� ÜF(��𛅂*"=�k���z�Z��֗�ko��=�/�m����,c���@jډꎄj���DJ]_OҲx�r�|l�YU������l=eܵ��X}_K��/F�#���I+��M�/۔W�->*��S�`�$_��d?GG����VQ���i�3T9����,�==�$Al�Y���'�h�$� 'Az�?��2#��ǝK�D�c6z~�m�fqn�ݕ�v�x �j�k+�������N���Ui���c�ܺ��� H�㜳^VM9Fߓ�M� 7s j�uA��/��֔F�Ʃc�x�YꆍQ�A����7a\e��x�hA~�`X�:`<����\R�=)��؉h�(�ඎԩLW�Q��E���Mj%��咮��:���
,�Ϥ��H ��Ľ{�o/�7�w\���[MChv.S��R��x� �M����~���z�5�z_�Q��rϓ���0i,�EzB��n�=[ ��n�\��CkՎ��0�U
�P��6r�3��re�1�EB�U��N][��Su
��uȢvueT���|�j>iZ�Y�KP���1�_p'���.vi}�8u�ʌ���O��?�*��ȍ��  ��"N�/_RESm��X��\��^�e{m�	�������\�ͦc���%��@Wn�g����e�b ��؂��/�x��N҈+����Z�g�Yh��9���T�
=p�ry�j���_k�UH��'��}{�J�&�Ū+}M��}ڎgd���Nr�.o��@�X����Vz(n���O�6�<�S�����|�b�gM�����;#j����ЬT5�*�NH�0~�<��n�g��v�P��~F��3FF���)u��&�0�Q��
��W�zgC �O�PɎxg;f Q�\V�4�>%�V��&�%ьPR���9܌��[)���)�.� s�k�l�\�J�� q��8+�{jF�2��i�� �ǹS�\�ms2�"�I�F�z1���\l?����}-�ݾ����wr�r^U��gJE��H�I�=��8�"�>2pC&�cI�U4m���������_L�έ�y��&sM0??Cf���<&`j�S�<#�U��0��M��Ӄ���v��!<=��f,�OlP�
dA9*��������ߌ�˨���.бj
��lAq�n|Xz�`�-���@��,��u��<�F�-7��߸�WK-�=���(v��+�W�"�ܲ�|6�n�&mݖ=jk^Ҹ�g
�F����&�P�ϛ�\O�9^��DI�Bn+1ī�����.)T�$K�wGǞ,�2�eB%��ds�����\�7AZ<��ԇ&�{��L�YwҿH��C�2h���P�	�g�Y+sU�f0�e�Y)nq�t
�� �&;X�6�lI��[k�8/��
�C|�������omM`��+���wYN�d�څ5�����7P�x~������1D[���"�Q�"@^-afH|��.���E�_���P�߅V|���T��	�o�ɸ����؟^]���V�y��|z�Q���h�%�j����T�7=���p�/��֢�̠���"�u�u]�ߢ�`b�h�c��H��>P�R�;>���?���]�u���B_����T�k��0"��� �4���`�t΍�0�A�c
��8�� ��i��p���܋��u9�	�G����?���S�y�z/����AK��g��+�DҸ+���b���<��*C���o����w���s88��m�Ĉ7
�NF_�%�`i6z����8���I�f�����~�Õ9CO��u����s��{�k�%1\)�4�U$hg��Pp�����X��Zi��~B�q�rJ�4"��*
n �6����\����?��p��F^�|�[oe�X���Y��Yp~�s�U�9����b"':��1�,)��)T��ti��X*ױC�]�q�c�05
;^lU����$�T�z +�ҝ@K�YI��|�/ � [0�R�<a����Cnҝ�ٕ5�X�ƾ��c���)	H�<z2�X
��%�����q�Xd���������.#B�Mb7bu�s���!���%p aPL�i%��0ʬ���B�� Xo9<�nR���l[j�d:\�%���m��(h	��&�f�Gn�0Ԭ�-�w��?��p�ڲy'KoY�4Y�ӻuvU�������26���vMu����x��
���z��u��A�C���Y9�,h��㩍{�� њ�\W�R�۟�����1�[i:�ї�R�P�$	��%��J��l��rw����y�|���R�g��)y聢����w�^��;��"���#F��Bƣ��ӑB�[�}V�����WFۼ�K�{l�_��#cFVD������F�4[֋-Q�Ϝ���qX8P��Yث��}<��#���'������<�z��A�HS�팲�4N������J&Ic��l
��ELp����/��:P#4W��#d�z����<���!Ő5q����Aԕ�a$����+���}@x�����E���:��l�V�?�F�A���	� Iw��WX�~dĚS�J�3z`�?k��n|��J��z�Q���#�FZ���~�Y.hv8��%����t����G|�9���3Q6��
���'GɟES=`�҂d񍥔�n��(�ब�.���H�$6I���uj��ڐ��y���z�\k=��e�IkS�XY��
�0NN�Cg��٥�����8���j��FGg�B<���|��rJK� ;b2�ha�.��&uĴ�߃�>�mO<�eK��K:����oj�։���Ih���冕�x���-S�]����$��m���1����Es���rI�ci���{xZ0��+:�`9%|7���yz� �1U����	���A��_;}�H{�wc��;#����rNhWl=`�5Y�o�B^|U�/w\�ȷ(�ald4>�S�t�᣺��[��QL|u�Sn�0}fVK��`:1L;L���	lY4$����g����H��D�����C��x��9��fO&?ڢK՗u��\J�US�mu9I������B���a�����-�+��b
v�qX�S�T��{5��
�hh����(���a��H�W�Q���p&΋��A�:�;�u�O]|�_i���.l9n[Չ+u:����n���T6hL��&����R��Bj�j����ED����8btJ� �xG��~�#��e�}؁HU{LQ%qw͖ �0�/�9]�7��ޕ�M��+�{x%/�92���>���;�aG�t��=NK/;T�P� ���oo��=AN��n��v�S}rP�q[q�=q9�r��/hZ��i�5aw����s�������@a��6 �> ٷ�m��.N5�b���q/����6����	�:�3��0M�J��$�+�I/ئ�O9������V ;)�}^*��QI��Fe=�Qh0U�Ѡ���8��D`�L`K1�h��m��c9�0���X��dU� .��9t�JInN�K�?9U�v�bT�,��N�j�E�@��y&֡�km���G�5��V�%���g��<�AFt�t
 =  ��Z�!3�P����T^t��B���P�G�I>�QhM؏�)J�ѳ�Q���Z߭:�&$M��i-��LX���Ɲ�Й:�Cܒv�_Ǽ���n2MCi�y7s I\G�_��L��F���~z�Z+���@x�4��]XX��):� U���B�;�t���##����$��IQ�t�
�Z��[�F[pH,i�5�0���23xz��F�������&����]�nقT�q�m���ׅn�a���C�T��َ�W�J������x��M��?�P�s/���F1���+uO�o �YJʋ��qt�\��Х9�%
v�j�����Zt�����B	��['�w���A���<]�WKF��X*d�6�|�G�O���`0����U÷���A56r/}�Nm/��T�/�ۗ�3{'��Hd��z	4�)אf���O=�7�b@ �C�;ME����5Z������x=��jbע���q8H�@��0�3v8�ް��Xc�;ņCD��F�!lQ�B�g��׉]�ߖ��3<��i]�=-�F���˰�s2ԏq���
�%���<O�g��w��>S�a���r��o<ׯ�$\������,�y����mE�g�38g���N�ӽ�$t�𢾻��/�r�Z�Fo��Ab<�<Lr�N�`��(�z;I��mb�	ϴ+�⿙�a��0'��N�$;���u��{ԉ�o/�
�u�f���'��K��c���9y�ȳc�M[��bh C�l�;U��E/l��"��� j=��'����8y�T$/��Ʃ�|o��K�@i)tK��OE�h�l:�NĤ�:��Jc��Lµ�\8��rc|LeKi�G��X�%���-���b�C����;�� �}U���V��r�ǯx��?C�9��Ϩ^^�r1g��&��KM�q�����Bb�VX1�Gr�a���ֺ�ٽ�q�1��u�P����,Kt�x���w�7
'���kπ��ژ�< ^j�Gec}��2���M��oF��ـ��e]���a}�Iٲ�[y�Rp��I�'}�`T{�\r[�ߖ�j���ȃ(��5��N*��V�C�y��Vx���L�`�̎Tf"�$B9
]ƊY�˕��O��*��=�c���H7G�����������
�+�&.C=��p-������G]S��^��"dtw��Y��������k�NsȓWK0"��(_�'f�6���i�t�$�e18 ��f Nw��봨�����3��o�ꔖc�&��4:��Ȗ��U��Ӓ:��D���R���H8?�f�6J�#��Y:�LI���^�k��>�]��:ŧ�̈�Sۣ
yO�w/s9�_��U�����Ȼ�����.���"��f�D��-�F7�H�G��d��|�_>b��2�YỈ.\A��h0zP&Х�+cR�Uݰ��A��lw�5A{�P�-�:��cHZ������'������x�v�kT�^h�@P`�4�h�����Xn'2�|p�u}��#D�w���	>%,s���ð+�t��"��"G��h����U���,����-����!>�]�I�c��5�S<�P0v���l��)�`!�jxZ-��#nƽВ,� "L}s�J����aṢJ=� �Yĺ�i2m��ҝ�W��5MnZ�U�n�R���'���_����R�LW��� �P����y?Sr|���p�	 ,B�w�[=�Q	]/qګ��R�	���2��e�j%�����KY���w�Mۍ����;����K�>���-h;&`��K��ΆxX���:p^=��p�{�ܼ��2�R��9t�G��lbpN|L�zeA*��m�~���e{W{IR)�Ѐ:l��	���T���v��N/��s`Tc�Q�K��F���r3�C�k��D���x��u�8�A�H��5{����*u�@�PV��<ۚ*#x8�R>=���i� �6�e��I��+u�+�����1��nhmP'�{9�]g��ø8L��/�wp��{�Fp������E�.>���E:�`��t@*��Y_��g#��2�o�f�ޙXk���9,���8��ѻM����E��<x)��S9��]ӓ<�J�1�i.6�	�H���B��NW��㪫��E͹_#l�������6j��SPi}��P��%�w�{��1sS���*�Zk��/�L��qM����!��i���Xjg�;�������& �P]0��9#K�SA����䁎l��1��m���,��@��4����s�싅ȘRhN#^���~��r/����i�B{#���Ǫ�᤬H��8� ���{������WE5����q|ͧh@eSȩK��MH�Ze�	$�j9"k@�զ���,�8Q�$����9�\1�{r�<"���ԓ��H?��:dsyS�2����m�FVӌ���R;�Wo�*�v4��&8���#0|�Ϙ$��b�Tq1QqjlC?�z�T0�(*7�����T����&�m�'xc&����C�5�S��hqD�����1�S4�VQ�U�L�n���oh�3��+3/z �"��Khn-�~\z�u���\�s�G,$���V_o����O31�B�䂱wϢ��PME�$Mנ�Z�w=>��G]q�Vꓗq/�g���ꥳp!���?v�:Y8T�H�k|�c��Y	;Z�E�#{$��*`��)�_A$� �P6��ndd�ϼw2 tҍZ�o�2s��Y5 u+�c؝��O��Q���}�mQ�n�)����^���9ߵ��/5�h�
>�	X/c�8����蠰��D��`�����>��Uc��6J��4����]��|g��o�d�1Y�j�Ό�W@T�ڂ���2��q	*�f�]��ŕ����2*�@ݥ82IB�Y�H#⮭�I��-djCK�"HP�`��!B
�:y�K
�˘^� ����B�kp�>�5�5̓ײF&�e��AP���t��ˣy���yKluE��Q��92xL�>�G�,�����q��$��">����H��m�<i/�nGQ�]�B�
�¸<��W�Qb������ned�
��� �HI	I{Q��4	s��K�d"Ѧ*��t+/[ ��Lv]0-a�Ez����	���V� �S�t��*�5�����
]i/+$ʧ����pE=gh���z���pr#&ڡ���9+��O�ع#��6�3ߖ��!��A���1�u�8�Tٺ�ν�b[��1�βCx�ph�_����_��i�����u �C���$����[�|�Ui#��!ԋ�H��F �d�op�5�<��+��13�G9>}!�%��(�y��m�S���,y��n ���|c�6}��6��I����WB�	s��+�u���/�<U�xb-3�G�ݚ�kq�d�ʪۇ� <�60�b��R-�r�k�g����b��3�ﯪ]٫�/�!m
�$p*��#�q=�F���ng�]W��y�M	e{,�\�>�UDh�W�;Ϙ��(e�y�X��O����S��}C.��zdx�~t��_�f�ś��!�U�
�X2�®-]3�sǜÏ�X�(׭-��ڍ�~�.(,�m��[��7����v��^X��62�����H*���1��n�(u��bJ�ш�xM�w@�O�"�0�M:�UEo�7�^� 5�8�H�������Q1��a^��9�N/��o}�sa�'DAs��݁2�A�B5��%ݕ
��� �e!�:jY�U�&Y�`0�<�P��a�｢����H2�пdT���֐m8�˅���gd��爧�j�gD:����c?֎��ƪ(��Z}p���,0t*o��JJ!#�� ��r#���.o�ǐi,���g�j��:�&�y��h�3���5� �SU��E�֫�g�?ŉw�{�B���x�m.9n���m3���\^��,�Н��-�t��1/F��p��g7$_���� ��������C���F��C�Ѭ��پ�l�WN�w�ǎ���0��I K\�K{�ɾwiB�j�(+�ھ�b����T���X-h�L�����k
N���r��s��ǈ��E@�V��z�٢`������Ohv}"aE�nI1%</@���4���?Fg"�ǁe��{U����?�
�o�u�uڒh��|�����o?��:qO3�2�[ɔ��#S$o�2n�D	tz&��$JEI8D�2f�L P� jY����x�E�/uc%q�`�J�;�Q8�G��*��r�����>��PQ�	y�=���+��#y�L!�[P���Z���4'�x��~̈m�Qw�h�`��x��ӕ���������;?i�u���\&��yX2��T�<h�ʚF�jepiH�&	;4@�Cƌ�*�3|	ߛ��SxgӠ�
�����H��/�F��(_\|�#���`^J��}^��?Ą_U�Ф�Pm�aa=��}UBhT;��ԉ0+�]
����L����J��g}����\�ڶ"R!Z�������
w�]�R��`2{�3۩�Xj�<��GgK���"·�RQޯ�<MQ��J�oX3r�8T���� \�-�lK몀��HlPH����rz��a��Ew!��b��2�$y�y�. {�E�:�'�r���b��J�З�
��q�(�n�%/����~�p#ᚒn���$��f �IMC1D�"�s�d,W8o������!d �$#�q���Gr�,W��q9!߁`��H�6tE6���i{駞/G����\j���J��<#˖�E.'���4 �Ul^ �FSp�����+���E�/�u��J2�)@�Z�����q+w)���_�~L��{�z"g�{�������#������-c���Vܟ~�C��HO��؝�w�b��2��4I=D��'�H��_��}���C]3�w<v�����b�
=�jG�R�v�pęl��������w2𚯎$v�o(I��f��t2a`�2�Tb�$�0D�;�C���'�Fq4U@���Y��v0@F1��7\��]���<�S�\��Ƚ�F��9������j�
A��sN<��#��}�4��l���5Hi r;;��4��9�@�:��-ôJWg{��Z̴� z9M�ѝ�˃�cU����)ͱ�G����+Y�7؈���h{��`1=Ѳ�κ>�B�7����X-�x����_�n�	|�tk�@�v�X��p,���1�n�=���������J����j/�,2Gx�'��W`,ȫT��w5}��[v� Q w���m�Ъ��;�N�oa�ƶJza���1i�p�f�1��w�\kې�FC�j$X*^}��}�{:��Xo	��ZͪĞ!�}N
Q��'�3y5;�$5�������t���?X@C3]����K�LU�s�0�?D9k5
�k�T�ƃ�aWHރ(��.�	I��T\�PY/�\ȕp7�q&;���@�TuJ?�L��7>���&!c�����"Ӹ��7DX�\�RS�۔]��d�3�u�wXϚ�)��v�eE��5ѹ��MI��E���n 	LP����lǺ��"��S˂w29B�
������#��\r^f�	&p�v4��ˍp������޼��HP�?�j��0|�_�l�/j�
*l�U!̡:�'"*3HvUƒ�La6�Z6\�@�`�ߩL�;�_Ѩ-)��smq�H=���s,��o�zJ��tm�C3؃���F��*xO�v��{N��e��������A��7VA#h�MK��Vݿ�&W�$3�0s�HOj����8����ci>Q&I5�G�'��<�O�ɪ�{��#��4����HL�th%�ֿOΚ$��ڈm��,�J؆~+��O�β��SR� �7m}�r}�id�TJ�v�BaH�����𸝫��.��5�sU�� 9����E�4$�(����=�%ԕ:NJ��izO, Ֆ1�<��7B�o�} �����(=����t3.�~�4������޲J�� -�tM�}�!�t�@/��Bl���*�r��Y���,����t�P���;e����~ω��2��
G�%��G���m6j�\��q���4bA�7�x����&f7y���|4���8�:��b/�������s��p�q٭� �y�L6�ʢw��/�hN.�Q~��Nh�R�*�Wp�Il���I5�PlR��O����p��6����-Q��ڪ�43�*��/7����)A^���i@%�����Ҫ�R�&V���3��}_� ��	"�\�o9���-$.ԍ���ߦ��m8a޶Љ&��h2��o-�cN���Έ�v4�<ӄ�56&���w?�o�H�P�3H�E٭Ӑ��4��}��&��pA�%���������#E�w����I�S����m �8��p��\P����6�����ҔQ�Aa�Q5{E����6,�*n.�Ў���w�+b�:s�aqjesa�HZ�ϫ"(3~��� ;$,� �W�z��.L��i��/�Eî�uR&4I�ݬ�S.e>d���i˵%ĪX36�_�����@~T���"�LW�d�y�JD�LX�.���i.]�x�lޔ�=^���/ut��r1�d!���+�F{�PDO;pl�{7��sq��f��y]�0�P͜q��n�$�g	VO]�/��_��c]%��wg���c�3��1-:�6���K��)�a�r�j��SW,���W��j�!���<�d����/���L�9��y�o��vt+�*C���.E?Oh����� ����q��,�b��ʠ���V�c�q	W8ʎ*�}ȹi����7�$��;3d+QrE�`r\�/����~�����뎪�E� ȃ�_֘~ �%�� ?
�"�[A�R���f�ܼ����ؔ����KF� �^R���r������Cz�ƴxL{��zr|i΃s(�Ejs�ア�h�D��N� fS��!�0y�·��;�{?�!._�a�n=��:�#�	��H�y��M����I�6[xݿ+I6�n`��7����Nhˤ�Ѹ��	k.�W[�q=�s3?р�׎ﭮ��V��vW��Ǣm�ܭ�7��־>_��������IvUP��K���a�E�"�{����s"m<��$/���4V�FWޜ.B|۪�h�NND�T6�]�^�#�s}�db��,����6�ߞɛj�/ܗ2G��ϔ��T�ٓ����E�X2�}�l[4��+*�\�əT�f���Qj�΃�%{��gZ`�#�8ֶ.$Z�ʇ|g��VB�����~��j W��iI�17x�0S��`y���zc�a�ب��h�K��IKC�gP?�x�i��s�Y} ��s�"Y��9fM ���������^����V��U���7��@,S��<���]Ec2��$�!d ��˾����^Qr��	ҡ'�h�;V��UD
�Q���ffW�z�F�U �������H+�`��8q/n�b�GT����͞�
M�sֶ*��(?=��*6C�n^g=�Aj@m1q�1K��-K��(�q��5�҉BA��FeRaS"�?�&S�Vܟ��>wQ���~���yE���悳7��7��)��@�r��C���_�� �B�"�LXx�A�9��([ױ�>�����]!o�,5��ZȘ�e���O��
@���� b��\*%�u1(j�*�6�n���H�z�߂c�,�d7�T>;�!�K{"�TԾ�]j���2u�?7E�*,Y��=f��Kq�����'�b���x��c�4�f�t��A�▷� 1\�h+�HZ3��/LX9g��fw(�U����Gkp:y<X�퓧����А��3Yi��1��q�Yö��~� \|��B��6s�s(����m��	�K�¾�w ��R�Ò��q��,~�������"9�@jڱ��!6�Fn�����u�)��Ď������t�P��"��3��I��'g+&�:���Q����5���񞏩[��£Fⳏ�LO��{�B��e������}�C,0���3�~v����	,�q�㺧V����#�Dq(�#ӯacHiy~�հ��¢���R�=C�a9X} D�ycl=J�g��^��P�G�y9뚫�x���w_a��SC{�"�0s�tM�ؖa6"s/�
�ַy��;�`�����zљ�B���t���T��@b�O붠0¤@M��ӼG�W�@�&8]8����;+R,l��A�OL�-��5�UXƌ�B�[�5�l�-�tfpocX1�6��Xx(�n_�-5Yfh���3�ȶ-�ӬK��4h��IL
�$���c�1>��_~�_��kE\Nb�ؒ
~C�
�������{�S[]�3��NQT�V���>�(�,Y��ps3e����
L_�P��f��ഄ�T+��G`�pS�"(4j�=��Vv�r	,Õ
N��KF~���� �+I4��|��R	2"Lj:	�.�	�����z��)��A�7eC	n�X7T&�Ɍ���j_pƲ��H3&{E����Sl���8��A��7������k�A�bm��)��0V\,��8gG�l}��8\�"B���:���Ӻ�a��x /��a|N	(����Ր���Z��&����X�͢��_���B#�������(��REj~Qt�&
�Z.X�����}/S�q�bÞ�Fw�]��!�2��x�6eǚ��k;5�mĵx��َ�8E��7\��X2Q�	I顗�?/J}+%ƿ���(W��=�qjV)=׽dyՂxoVo�2����AL%n�o�-����>�l����#dot`��$3�G���{�C�"�.87��$�'0+���!G��>D!=����L��O�o���f��n�tr� ܮЗRζ��!�hJa z�
���N��8 .�n����l�}��s�᳤[3�5/�Z,`�y����ϋS��5�#0'�3Ĵ�)@w�7|*����AP��?E�*$���<�����2sHֽ�b4Q��^-��?����=89
a�`Le�K�R%U�t@y@&��P�1�K|Y+Ȇ�`2�%]�PL&�,!�5Q�"�G&�V�A��vL؁#@*}(���eU9�FY%A	���-8T*nP1AX�=�gHM�K2��ELSZ,
s�Q?\������wT�� ��Kx `�i��+� �Ǎ:°amC����M�<�E��.���2�s�i���E�E��1�h�G�k:[�.ސʔ_�T9��
ԐG������E8�*�ӄ #	G��4eb:~h��QaɉD�����3ز#d�Ƅ�w��ˀ�����9E���]�l�IB��}a������_ݠå�����&�U�Zi�%���z�^:ٳ�	���F��?"��>a:�~ګ�s�����a� i����H�ߗy����F-��;6����.�{�j[ȡ�-$Ds�!���	�/KbI��
!A�g�r�46}�LJ�zV��dz>�H�#��p��Da�w��"�z쵌I�u��To����=nMs�󾮲U��%�x��<�ѧM�2'�!#2�U��e�y�Q@��=�4Ts�מ�t3��$P�/�kB��m��"����mU{�E�u*s�'�a�Of�*�]NԔ��K�/��Yd�[���iZ\�(��}�����p�+���3Zi.NȞ|��c#}ٜ�(?o�JF}��q0���u�O�ծ�[�s�h��(�����ٍ�ޤ�]Q8�A21�$sb��бkd7�(E�O����NI���`��,�:��
��-�Q����ֲ
���ww��u�>�7�F��i�.P=�<q��O{���۽"��rÆ��1�0�/�J�)�t�:!O1q���bb�����V��Fg ��|�w�2�cbf,���l ��w>�`���%�Ƙt���P��(�kcK
�tE:��BM-ژ�
W턻���D$�� �ۚ�	+��$$B<� �U�
��� 8�N�L��e�(����D���>����E!�_�z�!��?:ʐ�LEuP��p'OW�EU7�;�m	�ѓ���-��*�'�:y|��s�k��90��S�y?<�drSr�0��R<n�����`��:v4�'���Ä�d��L��چ�kz���Q���;P�!GY�r]r���S�.�Z̭O� y��C*�o��C��M�,%�k��c�ܔ:}C�a��{(*(�(:(���Nv>�puGk��ӯ�6K��z
PV����43v��q����3r)�L����9h|�\���~�St�o�:-֥����s��o�!J��E�Xk���� ���@�1tc����?��/������Q��
K�F%Q��"���ƾ+�i#�B�q�+˗O�v�\֎B1�AULR ڟ�d�hP�]��2�jy�De{t�P���╫�"���5��k��W|�OH^ʔD�cz�]q��ۻ�M���um9�]�'�B���9 ���(@⿾��[�vv7�a���N���.��-�o�'��{��r�]J7�gO�l�6�n�aD$�$�3n�
뀉�܅X ����{H�~	ϼ�jܜw���{�NƋ��6@W��}�R���?�\=�Q�b)��ډ��8͠���S*�>�D�*�#sr�����׾ƞĽ�,K6zY�`��O���hL��:ܧJÖ��RH�b��q�A��1n03�pO�!���Ȟ�QٮI�t�h���g/w)��%����>7���+��v8B�6ϻ����j��!Y�rmU0X���*��K�~�l�o�kT?u��#�W��zl����.,��4p̨#E+iRa7�0���>���0��D��,J�zO}���v;��,Lg�i���p�Q9���5ؕ��ߐA+�B=6�ܛap!X�ٽ�h,�]���M��u�_m�\�Pz9�0��3����6��|������I�Y̜��=v#<���E	B��>}o�!VqW�k���z|��;U��ґ*)�X� Jr�����=����M����q�>�ŷY/�Ǭa �r��7I2d���|�2�=���D��d�D��7Bl|X5��'|=J�y%<BWQQ�ֵ^��
cK���1`�+"�M�W-I+���"��$:�Ai	rn̸#_M'?c�F2���]S·�/Ub0v-L�ƀQ���x�c�!@�+	c��+H>��=5_�Qh�Y쮝�t?��|�W��e3mv�L��+�i�&ǎM�������	<�-NC�G�-&~��Og�x��E�܂?�FE`�ώ����k(JӖ�e�r_s�|��M��s�+�E
XҾ�,g��wC���mj� �0�b 6��!~d���6,ދqt��O�+���V���g�b���(�t�uݒ�\��/��-����ܣ�!&Q�] �姱�\��Yl���q�9�J;�(��V�s��݂\g?O�5�]ǵ�3kI�Q�Ww�lP��pI7<)���tCB�t!Ӡ�H��x�o$��v�O�Nf��_�Wl���q�Kܾ��\��fQ�Bx�ݔ��|����#�a)��*�gI�8�0�#�TXW��\],�{�,(o=�=��V&D���i�I�9�R_/���r��qs�.��~I�XP(�e�)����(f�������-yV��+�<"��>(S2�y���+Ep���˾�QZ[����䉻��@�&v
n���#'�+zz�-=�?7�I��[(|G��`zAe1������H���B�*��0�fĊ�G3N��<�㢲�����E�v��Q��%����O���YZ�}�y/�禢�����a �4����g�!�"�nk)��S��ꀇ�*F�4�_����-�-@B�}t�u�����9}�|�ygi���;�����ݑqEW{L�v.��PQ=���Þ��ĝ�Z,Ru��^li���I�фh*��apAn�I���i^~?�j��s���i׈BP�^��cΓ��CZ5Q�u/�#ن���ЭŬa�9G6(A�=w{۩_~ g���x�LR[؈5>��&MPO�w��Ǆ:utc2�����$t��X%?�W�}���¾����n(.����Ğ+f.
�9��@�(K�~{�8�9����`{�9@�e+`�4�ٍ �v���r��"�ʓ���P/��gճ�},��	�ff�22
��Bj��+'?��AD.2v`��UG�>�9��MA����8K�hW/���l�}�K�(z���U��r����n<%��cK0��g���5��W�|`���il���Ϟ:T6��a������v�!�E/�-3@��l�OG;�D:rJ�ț��S!� {�C�	~p�V�����`]A8�M�6*R.V��M8���.c!�e��#�SL{b>Z��0���JN/�������5o�G��Xcoj|�s"���y�et`�4< �6�� ��\�a&Q�J¤�k��5F��rbA!.	����)���:1������BI`�%[�����Ȑ���I�Q�+qb ���6x:�úf�K�$�D�s�!X��,%�7@Gެf��87���l'�U��V��V3�Yu�a���4�Gŭ>�!w*�d3�-=
���K�,�EJ�g��و����>n���q2I�4�$)�u���"�O�_�	=�5VU�8(a5��v]fI(�_=#���h�0�e�@�����,qfA�5\��,oR���=�\��U��iL@=�Q�.��h���[&�����������S7�#S#Q�k�3�TR�X��wGŅ�#��߉���:� �܀Nn���W���x�Ç_R�hm�9r:�`??߮Kmvs2C>�}����~pxvL=�s΍����q�8P���v��b��t�I��|�����D���fA�/��|9r�Oh˟}��;��EH�s�"v�������;��.�G�x�Md��8G>5.�k��!���s�"��H{9k����8��S����Y�.� kA�e�~Ɔ3��T]���ۮt��W���Mf˘�0O��O׶��t�z��Q/,2�H�I_�&W*���5�	���fi�x�/h�@�˚3����s���z�bۻ���P����l�".X��N��=o���'2(��đ�^0�rds�֧JtzV72Z�h�ˣ��GC�5ˢ����U蟓OYh���9��ݛ�e�U�4��⢁J�sD?���=r�(x���F��K{�N�y�4J/�,=��]� ���Yuf����
߄��S��]%�2d�*Ϝ�OUf4���cP9�5IK���4JJ����8���v�ɤ �T�cuR�-�Ɣ^ɇn"!�D���!�����Wksg�Kc�*�9TEy�ʸ+� U>_uP(�Of�7�L�������u禐��%%K�}6i��#Ҵ1�;8/�Q��Rp���~��5�}��xDFía���8�sC�j��{���L 5�E���5w�H�疋��1mx� �|����K��X�`� <�_��M��W�ȏ�55�t _�������n'��kFU�.�Yf���Vt��Nk�T��r@ұ����>��	 bů`��Ɨ�j/���m��V��ba��漯U��څ��VRB�|���t�UR�,���Oj^�av��B����f<�����ژ�� S���(�|�� z#��~�0�����kw%Y��N�q{'�Ȋ��K�k,�a(��RF,�"�k���1!�,A7ᑕ$2_ʦ�����y�����5�b�݇�X����ꔎ���J�����t
�e�)��cԚH��l�ܘܱ[��~	���_:�)�ɥ*�
�(I��1)��4���n��S���A�&�Q���o%��X��ٱ�mb}Qg�������4ٞ�"<A�mQ
"�A��L�W�8�Bh{y
�ôGP�.e^҈~�sW��^i��a�oR3�	�qk����׍
ᨲ�=��u$(�����^�y� C2;���;�;����.�S�!O���]Z��h�g����: �C��^��p��;��!���X�.Ћ�r�l8'^/���4�ھ�܍�J��u��B�h��=p��ZB�ƒ�C������xmoS�m���̣7�.|1*ж������D��Dy��L��G��O)M"����jhK	C��`s����b�O���\6$9�����vp��[�q����V{;����5&�%�,���A!�1��Fg�g��O��;�f�(���ZJ
��N�fP�J��[��Jh���i�gj�ˇ|F<H|k��
xT��4l��tG	�F�m����Hh���wܛ��~�u�Q�@U�ܪ#� ��U�&�zu��s��<w���<�QC��Xpo/����D'�M>�jyLطFt�0�I�2hy#�Vrjǻ�?�O��*|���~O�7��\�NYi�NK~�/��洨�;�Ǚz�'�%=��Ъ+)y��]���8��>����˗�c��"��Iא�����.�i+n���o/�����v��HQBn���eU'���|�j�fb��)x�|�I��Z������Ỻ�{|SGt��L�������uv��}>�7$Ӥ�D\��`	)�+�̍+@�y�Ng��}�C��g�65.T�=o�R�~��6>k�sr��������n2���D+���C���;��_0�'�7�G½�>�9�wݘ��<�`xz]���і[��$�I�)`=,�A=T�^ghJ�(��0��p�a�C���9�su�x�0r�wM���$@c��q�.t\��E�A=���]�)�8��\x��Y��u���e�+��`��oQ�MR�ֽ��*��ܶ����+��R�=�e[08��M�
Kn��+��-�*��<�ʤ���,��B���ؼ�t�{2� ��:fU��Oͯ�K�B^���~U_]�u��K[�����h�e���Q���r?N'��n�0UX��֟S����� ����"�����Uݙ�9����Y^�oW�=b���yo�7'>5%�'|g�V}��v�l������<�q�g�V<���KG���d�����st�ѐ���qd��2Vѐ���~���IYB��k>�̛�!!9�RV��;�E�E�(9.P̆'��ҟ3 ���T�9�e�϶�����F��"n^P]��d ��n�)�Q�:�g.�H*�a�p~Qp�ϚiJ�G��{�e��5� 2��#��9$����Y�ڀ$�CTl`c��T�y,k����~F��u�B^p,k�Y;�����Z-o�Y�Fiɶm�3gL1���: �eߑ��h�#`�&�,ISӬ�Z��"6�@Q�JZ���<&7ToQ
��y��C��爣���A��'��S�JZh_��]	'!�Mbu���^V�833��߆�^��QEE=�a�7Rcޱ��d��m��:��P}���i��i��ۈ�Z�d%o6�7PM����H�ۥ���=�\�j�����a�ǃYqG۩���fIC�=���ٺAO��4�)?�!�>Tv���á�5Lo$>��`�.��X�� ��?�Y�hp�W<O��6���b�mW�0B
�l�9�g+�>�aւ b�2�E���%�N�W��חP��9��%�p^}Ϡ�4D�X p�3�b�n��融	r���w'=�?^J�ĵ�%R�Ͳ�c$��a�c� :�(��#=$SS$�X �V�TNYo���Զ%mI�W`�}/�w@Ɍ����Ҍyy삃�Uo6�TlmX\^<���ü�*�"B�k�!Xc�����N�:��ʒ�1���Ji�y��aY���Vś�A��Kx�$'��,3���"��_�i:����}��W)���]���N�k�r^�3w��+������?,�f
w����4P�ˁ¼��W��$�ŎdJ��Å����q���Go�/��e<b�Wy}Me��jB�Í��B�PK��'���$
�z֑PJz�~[��4!6�)��2lav��[b�}�d*!EW��3����A+=�*�d��!䠈:��h �#y40���b��R��t���/Pr����W��f(�E;���q,�#*�{���sgt��愥�����~������!
��
�5t�Vp�6�l�|��!��q�C�,6(I��/D���$ ~�3m������������6�.�򂤰���J��7BG�S�?���������� �D@3:Wrϋ������-�${�0>��U��XםL�f��1�<|7��K���sM7\�<V>�,k�p��B��dN*6���8_;�l�D�H��]������2AT	�p<=��}G�ݐ�O��u����|�'�G��Oū�1�h��c���0�#n�!�$-��2�T�H7(/1�a�1RI#>��҈d��i~yk�0���߸*t3\$d�"�4(��>I2pn|�"�Ef:i�q��~W�c�$�)�����׌x�e�a"�vlB�yr_E��8F'~���>�v�C�JA���3jv�o��6:�e�|m^�������+TU��F"vMp��#6fǌ���R�<c�f���������OX�K�q�ӎ���lp��K���5�z��T�A���;�̿
JS-��#�NO�ƙ��p�KK��k�+�?_ErZ��(�Fn�)��w� �sr�<�/�}(�H�"����J�I��x
�2�EQ��%Ad�٥ee��j��Ŏp������f����#1AƎO��	������,�=�������܇���6�w�l�D�� ��X�
��K�3�w����o�m��
iF�\-��M���p{!��,Q �J��@3>�ְ ��`I�+x���bߛ�e� �}�+�֯"�ks�҉�����*�؟�̶��,��X������P~­���fJ�篤9���F�e�8V��������؆���`(���o�O��̻�����t�$�ֻ9ݾ� xph[J�� l�*O��U�6_��I@6���2��\d�7D��"0�s�j���to�z���a��в�� �4�vX�2Q˭F���T�q����S�+}��A3�����{�y5�H����؜&Ku�?�ٔ��Th�89�<��H8X�Q��+��<��o���ȉ��Z�`x�ԯ<��ϟg���H��5���Z6��*�6i�9r���0���.��z�2'���L�t^�ʚ��8Y�\<Kt$ٞT�������j,��H����t'<�u�Z��f��f=�oC�M�#~q���.��,��%�V3�e��F�&%C���D\�MӞc;��_�ٙ`,:���M�LͼP�z�q��`"�8���kk�v�Wt�N��ȡ���#1n�=\������\��^t
E�&��|j��>F��0`/�R	P��HY�@�@���j�kn�S[Y R��β$��[E���o"N"�ǆ<��M4�q��wNsƠ;�߰ss��^��F���膺l���KP5M_fv�A�@05�A]qL
K#ۙ�D��:B�N���;���m��q1��}uj����X��w�{;�C G�[s[��Jv����h��b1Q�MyX�ן��|�q��o��d����sU�IVh�˭�$f�p7�K���^�\��Ϧ���ۋI&�f�&�N0�z5�%����l�7M�nAt�-�pϹ2z�����xHUw���!�'$r29c(��G�	�#:�����!Ġj+#4.�ɭ�\��_��4{�>{L�Wə1���}r�R�k��g�h�fh���K>h�tc31t?) �l�����TNs������J�Y�~�v�FV�Y}G,u\;��3yq�B�pJPQ�[G���h���,?�2��:t���.U�+���iO�:�0L��E_����/��=���y�2�po�������L,���	ښ�b�3 ���
�-�G��Ȩ��ʛqe���Y��qֻ~�r(����)r)�oˬ��<U7&�u��]l?��[�{�ĳ���<ջ�����9_s`��#j��ò�Luk�8/SWN��T_<�'�e�r����ٍD��;/��CjR��a�a�R���߲��Tp~�p�% 
�Q�u�:�yU_������c�>�N3z@f�UZ�$$�ir<g��H��۱�$�~*���m����e�bV{��ɼ�zd�K`�'����T���e %w��RQ�;Fe�|_&h4���}��2�9�cW�.=r�F���9.�	�#�م���lt���#���Fl�t��;���ȝ��/� X� ۼ6�~m�rcF<�c�"�9�y?���AٌK,�'���f��ݖI箿�SGV���<#�E���o�מDQ�X�Z.��cM�a�f���A�L{"}<a�()
�B��p�e���uy]�#��-I�̧�?��B��;-e�q�'�0[���"[���n���W6?����Ky�b�� �m���PȼXm@nw���b�����S-� �!������Af�B��)��ns�Fu���Rc�oߖ��0����z�}��(�1Y�O������%=aa�v��^�9���-܇�ףcd�6z��=n"v�#���\M�k������};N*Z,p�(:sБ���*xbp� �X��3{�)Tx4z_�3	�� 疇N�>�����E�&>5Ȱy2h�����!h���G���*��E�8��Q1X0׆�9�r�I�v�Y�f�h����$I&�ɢ�:��ʭ@����@:��&h<&C?�����f�b�L�Y��P���w%硰���U�h���i֟'�b)��|#�d���-�-h��b��_5�
;��Z�(�^W�GI(e����4l�g���-�R�R�O-����lac(��=1$Fמ�,�/�`�	�r�H| 
uO�@�ң)Ϙ����Y�%�w�<
=����-�t����@@Ln����XjӘm�:V�3
�2*��a��:�J�^Lt�y� 0�����cV@$��d���	�B��f:6�~2^�(���"�G~^)̝9֦95�HI��¬Q��
�#� �a���1"j񶄬���@��kk��=�?C>sCS\�����d3����֋ho$��0"�o�$�GNf�*�O���^�%)zފ�&�;*� W�B)L�r��������]i�(.x�̄FѤ#H�a���V���A2��*;jC����M��Q�/�Q*���EǠ�j���}�<k�B�WO�^L�&�2��^ ~����� �5Di��&|X@{bg�4+�`�H�oY����E�Y��s����Z	śY�`j/��'u�+�vp�=f�xx���U;~�@�IB��ғ�>���'# ��y8��J -�~���X$��In~��3'�,�iԾќQi"��"⒪	��ᢝ��u�&>�a��x��`�OO�?~�k�Ͱ��Z7+��G϶��2���A�{p�X��s�-Z�R�پ���"D��z�O݆��ܱ����ؔ��V9/� �C^��/�ȸ�y,TY������g0��Yޥ �##�O]��I^�ڶQd�X4O5E��� 哪3UF-��G�\H�g��!��NA�{_�O��&'3���u�c��#D���Õ�CfE$���%|����[/u�P�h�hTXW�oWN�d��"�v�$���-��������];��jYVc��t��1N �*t��Y%��P9e�<��:�L���3��n����~���<��瞚��|Vo�$7����M�̽�%s�{�����<O�����E1<�KP�)?�V-܏N���dS���ƚPq
	tA.��!Å�������;m|�wt� ���I�m��=uA����<�H���9�	��ï���!�B����ߙ�b��ך'�!��4�����e��J6�I5'��R(-��lMNFy�y7��w�9��T��68���U��&njh8|��Q��*�	�3՚�����2�8��K��H���^�]ۊZ��a�V�H�W:��P�N��F�!q��Q��x��Y�0R�Dc29kh�F�gg8�:f/��)���x�(C����?7���ac��L�(�U��R������9�N�'�.ᇴ�N�$��
�1")ާ�ߤ\���~�]��>:-E�#���>�kI��ds�Ax$;t���7�˩h�Sm��SA =p��'�J����D�� O�����K����UD��-NZ7��2<�W�ih#r������l��Ɣ�{��O���$z},�Gf��]���S�������� 2��dA�Kބ��h����z6����>�"o�K�^�B�׮�I���oWSg�2~V@��y�,�$Yד^v61�ɸ31�X`A#c����r�:{:�M�l�ݘtJr_t������S���5@�@ˏ;�p��B< l�0U�!�u!�I��
��=���H8��F�!/��k�q^��e�7�Z;�=iO�P�/p�z�~2��R��M^G�������9z���y͠����=���~�Wv���5��D�0�=�5L��@�2��dwγ��/�X�*Ф�Ag��q@m�oE��H)&P�.y����!�#��������u)��(��Tՙ[���~x=eV����1̙� uӒ{Ҽ�h�zL�����_�q9ш���p&�f�<V�����h�+W�����_C.=���d��e���d�{Z&�h�g����.�.�T4��-�O�=V͂�+��� ����$�m�de�(�WD�Y��<G���:$���S�\���U>���؅'�i�F�=�F!+/��@K4
}�.�p���`"�P�0q&��3�9�['X>��C��k	Jidހ�{�����z�W&�y^=>C_'0i�po��+S�Ik4ٮ>{LV��x���R���5��ͻ="�7ܐ*`�2�c�Wl��J~.�(��f�O�/$�0�|�sSx�G�� ���G�h�议�h����bAB�ŭ���L����BV�����ʖ��qc-¡�++�'��:#�b�a��S�7�U�ҍ#�Eѕ�K�@Mg*2����.0 ���඿��!jH��"ט�����6�ơ+n�q��YE�H���ym�1�K����v�l������4�U��+=�>�]����',��?��D%�*Kpm�B"�M�]Y���D,�M���pA5�i��>/�E���q��(���xY��ܳ�����#���/I�����5��RIR��=FY7v���q�+\%eK?SDw��gnc6�u���g֫�_��I������a����NVU��;SZ�kE���V��J��;��`�WV����7~$v���[�Ƹ ���C���b4~�����C��+]�eE�m8/lw��P����Й�������7jh=q��M�
{�S�)�63��u���+NN��ƨ2?��/��/ܟp��x��-k�Mo�}^e�qvy-�3B~�I�	��W��Ik��if1���t���4j��wi���tBv�~��'�`���I����to00]����6���&~�vx!6'�c�~��Gk�(<P�ͮ��e0����@\�?ޛ�8��.�%�q|eb��|���������p��C�}'�|}Q��ep0��>�W�@D@3�2�ψ�\����ڡ(��g�d�������U��E0|����`��*��+����'ʡ�h.Z��z�jR�Y��g����a���뇖�}�YH�W;��!���W"ĝ''Ke��y mJc�9M��������1>QCV�)��6d�Wx�l.�-X����Ƶo5��e\���o~+2Hnӹ<
)1O�m=t����^G��:*��m/!����~�`� P��W�׏)��?>|^x��N�6Uc�����H%?,��7������7����q�)�&�j����<-$;�E\��xT�̧�L���;�wL��?���ҟ��i�pA~^G��#o �-;���@�)\�ʊ���&�wAA��
I��A�p����J�y��Pћ/9�_uY l���z�N�Q2�Χ;~-�`�% gN#~��֮���� ��5i<SJ�>�ΘD��oDԄe><;�̠Ϯ�`W�J�T�vK<��W�$c���T�q~Vsy.��akl�����C䱁�O��.�H�[�g-���w0�L�����p$0B�S�7�7�B�u��t���:�eu�;�o)]汨��!��w����몡}�fH���
�[�*�8?~����@6�9?yD�Ek�"�����P �'��P�#Wc��vT���\HtKYr��lU�B Ea25:�lr��s�	TQw0bE�I�����|o�m�W`j8��{�"��G�[*q�X��)oo!�v���[�+g[�x0(y�����W�M�Ҷ>�.W��3��f\[�|�L�p�J�V H%�C��W$YO
��d�?|:c��-����X^�~f����bBA�]�{BS������ĸ(��my�P@�}W������xh���[w,���\V��K�5���9�9��^�(��Գ�,���܂��(ʦc�:���hR�_G`�4&��� �AD��ɧ�Kn5���,6�v�G�sm������E��h�pbX�V�v��%�5��wA��x�}�|���C��EF��uW��Q�K�VHu��gԞ���p��ɉ�IV�pt�S�le����3�_�+O����е����&ڰ��ܕ�6�#�;�?�oz�"��"$Г��+b���
#��(;!S�u��d�0��U������ųSy�ᮨC. 5��N�d@)���W�CMht9mW�%��n2;�<Cv�#�� ]�~�G��ZD��ڭ���{8
z���e��Z�R.}�F��콪c=�6���c���W��j�N��;Dmg�ND��J�v�o�n:�Oz���鏣��V�Y�H^霙�*2C�,~��|���`۩���/�{J�B��t2��6��df����M-��`^�]f��[��ɜ	<���_��[O.�W�Y	��~�&�.2n��Q{H�1���
3kn��1�%%�1{O�?6v�f�w]8pW��2������	��D����B%0�k�kD?*^�U���t�������J�y�㈣��&H�	�����1�s��V���.dp�R!��r! j&����p�Jo�G���hr�p,���/���+��Y�6�|�f!�zC��~�,_���Hc�]�mM�� ׭��˃Cabn� �q��XqzXz���1���/�XA�"�F;\�$�7G��SJ�Cc�"���G��)u[O�-���k���i_�c�.�*#�#�"��PO���W�O��ߚ��p�Ǌ=���!<s���'Zw�W�-�Y;�������x.e]��~qL���dn3��@�I&qF�o��D��Ԓg��Ӻ�~����<d~��Ǐ�IELک�'� _/��D;�}J��a䧸&�NOU�p'�lD�� �>+��U"�䅟�83J=x�[HF@�H^��}E���	�|yG��']KJ�S,
f��J@��R�Љ'�����A~�@S�@?�l�)��*�V�P=a�(;���@cM�mM���"Τ�jՑ�0� .%��}�d�x�=x6w�7vsG�ħ���>ՠئߛ�79]�LH�H�	�^�M���j�I�}НS�oE62@8YrK+�d��V�]ƞ/ʃ�[�x�N�fZ��Ϳ$���(`(Qa���@���7�wm$_dx�@�_zΠ��Ri�πK�B��ٝ�P�y�D�'/CTR� �^��XN���ܿ���K	uM��ϰ������J�	Z���z� ���C1�A��±X߃�.gZ��u���HЈ�qS�'��G�Q-M��n��e1��B��
a�rK��(���V�3V��*���(S��^|@r0��"8����w�q�>��y���.}������؞�a����y��S�n��
��*T|�/晭+�ɒ�H(�*.���rsU�%%�L�+�J�N��ؐ(|H����o.�������G�­�vG2vk��p��=���A�,1�++�a'��������+$v�P��"Xz(:<`u�V��6F��{���	�onG�T��q�y)b�\^��$��pb�{�3A�'����׆��r�k��Ծ
)�,�ӫ��`�o����+T��� S���}s�/aB㻧	��U�k��#:�62�~�_�_`(0���H�g4c��ڱ�}����V$����� �[��*��*݃�#x8��2�m��^A�a���R>^|��9b�O�w��VK�W�֞�+$���!��� U,�8���\ٌ�*Y���5�o#;A~�^x�}�c�;�v����,��q�V�k�Yj?�m�����"$VUSX$�YG��{�~�a9,$7�U����5,>��zT��wjߌ����0p�M���g��J>�d�?�����4>�~�ei�ث���kF��^�K�����w�"�Gg?�*��=:xv?d�`j��k�=��iQ�f2��W��3����$���@�oG���Tŭ���0I���{T5چb��(��f+�촛�0E-��fl��f(fmN?�J��"�_-goCP�`8�����+��E�m�+�(�#o��k��|��5z�_o)�0��pn<Yu�[�	0��#���%kװ+ןy����GB��}�ٍ�G��M�+��H��7n:�cʟ���s��� x��:�v�V��[�n����dRZ���P�ǟ�}\����N����N'��^�2�g���<�O*����yP�w�����	v�h�Q�j�NK�����U��7g3�F���s��@�6�8׀?U>ݦj���:��B�7�z)�Gh,�i�����u�B���ek��_�����<Ġ��s�<[=M�ńf%���Yr�V��}i��C�#j��{ő^{=б��ۄ<j�I��A���\W���x.'JT2Ƨ��S�N�m���p�M�nwas{YJ2���.B\�002����;/�a�WQ�U�����i��u��G�=��x��Ra���4@�EZ㧗��[=
۟���+VC����s����G����7{�PS+�@���E}YQ.XN��<y�}�����h�!Xo?�u�M���	<�Rl�"�$7���P��>YAg,��}��!or�m׉��r3F��·����}C5V�q�0)p����SeL�\���0A�7��	5�3�R�l��\�W�3`�E���P閄��	8�_M�v�t`#N�MԆ;���C������놬���D��;z8t@ڈ9j���c�쥛�\����{D�P_Ҿ��r�+t��R�:�m�./ridN!<uc����~��Mܷ��b�����u3$Ŕ�-�����;;7��E��Ȅ�G��S��B]�p$lX��� r ڜ���s��j���@.,�.��2x���&��&��x����u��SA�m����Z�&W���3��-�X�4`VEN2�Dz�ˉt�,B���*�'���U{��4ѱ]��PE|ީ�)�`��H�H��NA��������\Yp�o�q_�	^Q�ɨ��\`k�ё$��ړﱍ���lV�6��8R�9��g� �c"q��$�u�4j*U���7bhiZ��h0��'Z{CKI����W���`�Y^���H�<�R���ĉtF�oϤ�[G7���L)�����?k���6�[�2X���8x�6~�;�:��Uo�M���J?]9� ���<��%�9�6��ُT�3���`��e�� �8�H�]��@"�DP�5+@'�8�$�Hot��l�fד<%v^��6�����>W	�osֻM�~XA���Ws�gYG�~�t���Z�>(�h@J�u^��R��֑X'��5�ZV���}區������<\R��S/N.Zl��@	Q�����HS@'��{�R�JY����S��]ai�W���:�et�� �Oz���l�?�s���w�}l�6�M������!w�.����N�)]j�)�@L�B�}VnN���3�h�ؒ���qڄjQ\�|.(�:Ɏ7�G�XM��2�����{)�@s�|n�ǯ�R6� ��]�����)䡽FyFp�����#@8�o��|�|g�a1�8�_c�FW^Z6֒��gP}4׵�g�J=߃��[l0.B���fT�J<d"��uYȡ�_[ȳ
�l���=hhɈ�4����AA{�6��n����w����BtWi�~����&��g%�����1�eA� 9�b��3�x�[����xRc���(qi��,��aC�v�C��6�� �"�����oXn��9�mHE�V�e�G?ԩ,/�Rn��>���4���>�%T�D}���rF:Q��c{N��kbzK{���G���E8��i���i��-��޸�y��Au|ɔ���)��4{��m9u��w�d�I��i_"���]�O!Tu������@+L��V��>���gnʊ�+
�E�LI�4�o��ׅ�m�+?�`FJ[I��.�W<H�U������@����M�@b�P��
]�r��Ŀ�]&�u�T����Ф!蝺$^R*>�c�du�$̷���*��կ�&���ڻx�1\������Wt5�xD�".�߮ ���cc�P��zPm�8��FtCI�}b\�¼�Y�Ƕ�>MY/ɀ�Q�KX�T�<~d�L�ب�=v����vħoנ|E$��\7n�|��Y�Ҭ���m�x=�<�C yxc��7���?��A����c�vˋ��Hz����w�`�3GQ6l_��ރ�k��S��Ǚ��p� �r����`�������3]BZ�@~R�۱�� �Q��5�-�E�.�a2���� ���_
	^q{T�S�8A1��_���X8��vn�|�'�>�B����t}�+��~���Ta)��(��;P��ș�ZZ����"A��:P�v2d���1w`+����!Ϸ�9��o-2!	+o@=8�����$�.�6��c����.�<�OZ8�Fɥ^�xaӸr�Ó�Oe����h��-� 075�lf�Z�<�s�Z���J�jkq���Vn���w~[�_����w��0���S�O��rſS���F� �]c%�������;@1�r^�%& �(�d���E>u�9S�⺁_����|J���|�%�xϠ	�}�2�����6.Q���b�Og�km\*W��N���X�X&���<�5��З�;�F�����@��W$K]d�7;�Rj �l�s�hC/�غ\��*�Wk��J<�y?��(�l#<n�{�*��DA[Z oP�`;� ��I(i�����&��^{�INƪ>�ޚ�1Α_���i���YVu�7�sj�,g�u���ʶ�y�q'D�a�-�a,�w$
 �� �"��]ѨŚ��������&e���ʂd�ge�nҋ�[�~/�ټ�X�"�-��([��J���f#���&7ȰS�'Ӈ����k?�f�Wǳ�/	9���Xk[?����V��� 0f �-	R��FC>��yD�y�r�6��7�i�;���v��p~��t2����F��D-��rϐK;a��.��}���3�w����"���(���3�<�~� �� ���P��)@�[ϩ7��V������Ϝ����"h �%��W�8�d��_,��d�4�ٖKfWw'J����@��Wן�f���VC����c���1��';EF��v56��,�3ήԋՋJPZ�y`��������mj\���͡|�p�鎉�>|��sVz���_k`�����1�_�L�0;������q����vk��CŽ���J�M|E����c�J�m��$�-�'����pE�[�*��&b�9���8�sM��vpK�>���&-���{Z�F��v$�L[�x����~�s���ж�c�MU��7��+�gˀ/�O�ʥx��	,8�]͍?�3�������_/�i�~ɋ�(	�Uz�P��dЌ�j���1ċ��C\�/RYJ��q��E���]�J��q��hN�k}�+�����[g �J��"�N{�Q��h�{��)r���ϰ$/.d^k��*RkS�QN�����_$*$?�HW{���mXAR6��\��m�� zH�*ĩOK�*��F��Z 0�w[Eu�>KBy��e{��ޥS��[��0�C[��e^]bb�P(��/w��ȃ�����k��&&��C:�kNjQg��U�x�� ܙ ��I5Y��	C�P�B��z��S�ZNy]��@v�i���&s���nregCs�D/<�y�Ⱦ�zf�BG�/�s]��PQr����'�3�2�B�l6��H!b𕔣-��/�Kk��A�U���$t�������`'�T�v��CΕ���).{7]؟�b�3�F��H�$d���*%����J9J�6���J�;J:���+���=��>֬N� ����MQ����ZW*S�����:P�������ؼ ��˓�:�W��}~h͵����2�E��w��S~�]g]be;��u��w�n��5�`�2��� vErX�{ɞ�낯�@E"(vR�_6|h'ְ��_[Bh��:#�	�	�����dk��L}�ާm�	_��.���'����A�X��͖��E�<�ԝ���8�[`�/-D��RF����KٰD^���h��us���ڴy����|��Yo<���|�o�=��w��c3꧞�_�<�v~lu'Q�2�Gy(5Q�,Q~߼��dX���=��(�ػWSM�$z��ԴR���B�ɮy
>wB�b��l��\ϥ4?�|o:#)�� ���Q�a���8Z�5.�m?@�⋌T����B��1{uyNy����D��'���C(�d������T�]/�fO�w���Ƌ+9���J�My�Da����^�ԃ�8�a�5p���ev9A�%%�Uf�G���ݞSo��KthA�<n�)|��,3u�(hO�]�D�E@^^.?]V���X�	��`%�ie��1��~�V��!��iߪ��64Z�W"�"kjG]U����r�Y��&��:>�7�{4?���I@�`	�O�W�</��64R�
^�����)|�"�wv	�J�/��&��}q�U����тN����F���JS����^����K_����7�E��xu�۲Z�ؤ��^��8	2,C������7m�Ú�6��[d�eP��7(�.L�������R��ַԎg�_���Ho�oZS�/�U@��b����o����C�,��: ��O�xe��<>��鏕��$���q�gv�qu/Ox���m��qth�o�2W�{<�(s��Eh��{[��҈J}q�5���%�K�$95b�ғmV��=|/+�l7ǎa;3!'Y��5�{`1Q��,CƿS�����]C�P�������j�tM�*�ګ�1��w��*�*aFTjKt����1]�I�)|@,��,��J6��H*8�Y���� ��(���k�m,�c6�=��$�Ld�|�]5�������V��x��&��*��ڝ����?x(Ƨ�*����^�*���~��zgі�ℤ��R6jnDc�n�FD)�3/y���eZ?&����$�mM�rpY7볳J��5oV\�Vy��h�bEG}�I���2��=� �ʨ��[���tT���rq��W¥�p��b\��*	��&U�	{�uZ����5�o�S$݊�Fף����v��>�ٲ+_���F��x|>����B	+��HI4�<,�Q�.,�&8AY6h��%w��P���n��tNjP��v ����y˱m�mMfۇ�^ ���>Uk��]��!��t�)��c�{(�o�	�+�Yځ�f���T���g|��Wڐ+3?�}n��PѲ�W*c�9v*@H`���*)ֈz͑��O����r\�Xz���@�����t$;�w?�� �H�'�x�,?��9�ht�̹!�`�R����+��u�2~*�[[�CHR�Ɂg�A>��EY��=ix�Ҁ��A'a���W�\f���C@R���E�
vV����tn�x���"��x5k���I�.d��l��t$��#�(��
	@�F��ߵ<"���M�2{vFD�+�x~5~^��(�@��R��,�S��#1�}q@V+`�g,�QQB��z�H43�'��3eb�ȵ4��f�p�C�Z\oM>�.w,��|{p�Dp�@����Ж�3����`J����XX�6VV���昿̢ᢋOā������<*=0�K�A���r�$���Ѓ�v;r�	�)ڃ�N��ӄ�1�B�fi,��H_�����"(l8��|pձR�m@�i*@��q!q�y��_�l�����f���L�V��rg��\�q'���N�3-��.�ܻV�S�����1��@�\���[%�2
Q���϶BA�\N4������%+�U���u1y����ݗ���P�}Z���"�q
�״j��5P��!��B��ʗ�K�I��>����@�^�l�٥�eC�u+�t�}�pU�okX<\;�,�nD�V��d4� H;!����^�U�bu�5;c(�4��4�٬�=N��$pD��g�u6�K�(��͍�wr�����zn����_��o�������v�$���WЯ��4�?�N�U���7����(p�e�P�����������@N.������H9�^2U��)�$)������� �|���,����*A}��6�>���iGu���.R���R"h��֧t��Ӳ(��E\�r�Yt�G�d|� |��Rh(���lN��&c�.��W�ӊG��CM�����/�f#��[�{���DWN:4b$��{0}���	��V)�H�T�e_̜�"����D�F�l�4�'0�F�~mo�����;J�K���:�D�Ē���f�ޛ����nu�, ������!˪mF������?c+i�	^�>�}��뿿� ѯ�1�S�b��Oxl^� �܅�+4W� 7��T���7�T�>'*%��o̤��_�)�G����b������ӽl0`+�\��&r��	+�t&NK�f4�$fHxC�8����x�������&���=1���qb����v(NC���r1���b^n	��I;X[���SvYJ�1#n�tC��Z��Z����w�9F��D�1Ĥu�D���9?��T ͭ������>e`�Ns�F|��_�ބi�b��M��LH�y~�K�x}j�P,��)e;8�U��Kp�i`~+��o�`�BS;v�Vc���4zt^�Ũ�z��^ٖs���t�`��>=8��dڠ�'�Т2��n��2`�Mk'�
�����u{����x�qgP�$D��ܕ䢬����n�&���74�TN9�x2�+��/��k��s�nV���[���+#U2$8�l����u*j-Li�p�9*��UUV�7yC���xN������h��#�}�1�o(4I�;�s�3�'����U]m�Ld���NN�}�0����P R�X���^=�U~p�'�x��>��O��U{��%��(r�������ܲW�X���q��q��ZtW�1�����|�����^�1�.��7I���T0��#좩���3�^(�(�ߙ�$�B�l�m����@M�ic�r"X��%�i��eL�q`	�d2_?јW�k������sܑ�]�p��X{�޲�Oɏ,�_���ي�LHu���3�I0�h���������b�,��K
A!X�gEU+TU���v4����X�C��ZuX��FF)�B �g_q��ǖ�h�}v�&��g����R+��^�¬�y�/�/�/;��3���%�i��=ZF?e��!w��G<�	���m,�"�B~��~�IC:�S?]����|W*���ه^�5����!f��鮵W�U�Tm�9�yA�0b�ϧ]��|$��o�ytS%|%5����ܖ������xvj��d��,�H��3.9�\��
�;.� ͝p�wa�[
�/Y�^��c��t��+h��X~O��Nfâ��4��; �[�d�|*CYekw��4h0�?���>V#K��;C9(�X�>����C���f��
z���W��#
�����v7�pf�"���0}�aUD�Z��\U��I�H�Ծ�QB�L��G�%8�v��I)u8���M����f�m94[XL����[4�W)2혼f�E��P�{c�3�D���u���z���#�%���8�Ѷ����z�Ztt�q�.��*/�sХ����D��\J��,�G�N�s�VhA�6}�Xa��+�*���O������"E�b����HK���C�v�;�X�s���c���%��};�Κi_Z x5���_bG������7?�����A�0�������?�V�C���=���(�y�?�V��D��x;6P4����(�[~4�xӅ�2��@��T6 O��ְ������ǟ�l8{kU�:�x�?�����HD��WMˊ�[`�46š��+L��rR�R����������WaךeK(Ʉ1�4��$.zM����f�5�'�r������M��$f����nb�箣��khVv���V��1�~�\5ݖ-Y�����uW�#���Wi�,�խ
QS[a���G&����	��VJ�1Flp)49-L
9��v��$%c���� fTV���ZG45���D�D���@��˲�`�G���R//-&��y���Q?Ƈ�z�7�z�ͤ*x�UHPZ��5e�����a����������2&�#��K�	k7�9��v����Am��%R�(p5�l�����V���%K�H��O>�(��ň3F�{��sT�;���_}O�原�]^�Z��r�Ǌ�������k���ߢgؑ����� =�|>)���l�y��U= +Ίܣd�z7A����7A�V�h>yP�Z���ޫ8�QXgY�i�#N�b��|�����&M��Mݳ�~�j]VNV���~�� �ت	ۍ����3�a�q��\s��&#�5���R$;��	�9=������ͳc�7�Ϲ�=*`�}H#d��5H��0�x�S�+���,���9�^�'���z����9��X�n5�>b4y���=2��ݢ�-k������1�],<.�N����
�̗Q/����Ȱ>6�C��� �t{��(�Q�G�+�_Ƨ�6�Bvᮠ~��;���^oa���i�����m�9�	���m���Ϣ���o��Х����C�ڣ�j=�4��rV.��ԣ;vN��Oq�f��FqN�	��&n3o��XHg$F�%e�q�'��_4����]��dr(g����X��GA��ܕ��[̯����-�W���;��rռ�z�ʈ�3��m���Ô�v���<�3T^�D
��\��=�� ;7�����!�u<��CV��Z����Z���ܰ];�Ir�����8ud�a\��ɩ̱���#�Nq���~^�b5L���C��`f(�6��׌d��[`.��N��˵�v��Ǿ�6b<'�Ug�n��hs��!��*�	�m����.�����Xnr4�}�T�,���D��)MAA���"���CvX�����eV	F��73}��p��7��0A�8���&�
'r�N��Cqn�������D~k���
@�#� nˌK>Ɯ�Dy�rW�E!�̈́�`��MP�r�W0�d���C�wKZ�3aBk/�iry�k_����]�$\�?s�4E+|�W�ɋ����{�}�(�p0�O�MAX�%��K��pD�zʱJ�2�D�e�EͽOK�����3�wJ�~��v��媟9����V��ĝ��NZ��2�v��͊?�hSQ���r�����$�_���%l�I��`��x��-X�U��*�Z�!��q<?�Dq����C	��d,��;PB7Y����OM4��*�����̝��6�ъB�6�?	�m�����}�Hs�Q�'��@x�=H�!G�7��ٓ��[�]q�D���<�rX��Z]G���%���D���֍��|�)�vc���M$���K��1/I��[��V-R<�l�z!�"��5���Z�tn$ �
�����dTN ��&5e�v"Ţ�M�},W;��ÐӨ��"pI��y�sGZ����FQ�l�r�s��{��K/s4����>� 䡈׽�4��Q��0�lc�o�i��K�^ ���f�3���YJݫH#��kc����4.�X%/G�k|8�ԙc̄`Q�p���|"�i-䖶�<:5�?���ӆ�$��a���;`=3�{X]f0�=ёa1��zz-x��gZ��t���s[�tRM����Jw����Q[!���?#,B#Dc���jP���^��L�.�8���,<��fQQ^F��� �6���-��z��
������qQ�P�=�8P�r�P&�|mMA��A�z,H���8�����/����bqw{K,^F����@P��~δJ��;�����.ۮ���k��y�]�8/���,�\	+9i�Dm�21
k�D�دt.Fez��Ήm?m鷮rRK�Yj.� -�:��t���3��@�� �^G�����K����𘬥� pA�h:w��R����%o��[�pA�+Dy~W�NLJ{�S�Z���Ķ�'R<���zC��e����)f���8���J,�:#��Otp-�mu��C�HV�7��-��w�]=p厀�3 ����}��	��͆���@b��`uJ���e�t͋j��3��L�?��X@Mq*g2Ƌ*�M��E���:��P��V;���eГ��F��=���mƷ9+�>��yc�-y�}�v�˔�o��\&��ŕ���I:OS���>U@���� ���h؁bzk��P���0C��=f��<�/���%��͊Ps�� vk@{�������FU?�,��E_�fw-��H�M:���0֋=���ʘˋ�{���Q�އp G��.C�?��~���H�@϶82�{�R��Xښ��g�f�	~?�"7��]4��&���+Ӻ" �{�
�DGb_ȳ�֌2睠*�ڀv)0��eU�4�w�=�}�$F�35(�-$V" Qk&B�bV��c��_�Vֶ����~3���*J���U��T�"�lw>��|+��T��W���:&�_��<��A,�b��T�~��G=xe�b��OD��o]³"��:m|ġ]|-/��t?K�IC�@�vP�&�n�����l��❸���h��m|x2%9��f_2���p�.�ڹjy���w8[��[�6�)&f��2�����4ڎV�iJ����)1�po(�����׽\���B�h�? ($��WkX���R��B�P�~G,�5*a=q�\�n������v�L��a�x�hn���q(I���Nc�L�$�H�ջv��d�ZL��s�x�V��`�=s��!*I�Iw'��b��[�s�.fYI��Z�a�A�|-�d��zkQ����@��5�<k�4��	�~<�+5K)����3OC�o?��!cO��5!� |?� ņ�37]^�ł� 1k0�J�f���ʝ-b/��Lr��-�4�H�i��_�-�r�z�]���Ǐ|� �7�����պ��۱���Y��G���hn�Q:]��-�:�=�)<�}��̎F��D�ŕ��
�����ty���$����襌%�\���&V����llP�R�!p�jy��x�|G�U=�j� 8��콹;��Kث4'�vP�sve��s8X!d����h��n��R��-&��=JO�HLBݼ@�v&�����p{@5:�έ7`6�JD�5tWO`\�B��h��� f�D��c:${��B;���;�t��6��k�;�a� D&����{�hp��ֲMK"�͵ޒ9���;���rw����-�4�$�Ă�{3|������t��m�P�'7�m�#��L��W#�GǮv��&�������֮UK�l���7:C��}�GV�~/4�@�,B��5; ������F=��֗���"�	�e�`���\�LS�8i^f=SE���G�6�!-���S�6���\���H�ȉŬOÝI�~��'�M��	�Uc	�
$knJ�Wǽ�m����9AH�`�pP����N^����Z+�Y�_r��-`U�����aq.�݇�#������p�n��/#��"�~N���&��[�����i��$�����aO�!������M�(8�q�'�
u</�B���� �_-e��F�O+�[�|~a	�(�����ц�M�$��^�>���$�[�+�5��6ϼxI95)5��9�tD��D9����XZa�e��WA8�ؙ/	n�y %��B�'�n�S%0/ߠ��/��U��]8�㠱�_�?(f��Ho��֩݀�"Gu��i[��F]�?"�k�0,�NI�E���+��[�Qn�vn'@�)����Ȏ��3.�1�,���d�w#$��5XN�L��B*>y���'�d%jMݞٷ�0���0!Y�r[s�f�D'�q�h@X���5wf"��E/TL��N����-���	IPL��ʟ� �Z���@�����̟�Y�����\�𔍙:�?�+��>��e(?8��{[�}v�&�`1�>�Ԕ��7��}��-�r�v�,G�6j�j�H�g~w�Qv��P����s����hI��n�=C|jo��t.������.kd`�e]��j^�I+\�x����o��� �R	^���J���M���q��
��m�=��:���U���{`�T���6uB���7�5�dI۶\�k�ǡ�*������{�$��5�L�/F�6k0�6�V����Vii�H�.;<�a�m/���/'�x���	
��Xs=��}���E�n�zv�T�KI(�'.��"1�(H7D�@��2vJ4N.��+q���*��;nD�X�B�hQ�%"�����
4�9x����g$��E�*�`��`h�q�a��g���8�P>�	��7鳔��q{N�(�nT�vO�{��P�]E�;�)�;A��Q.�9g�$��T��_��[���6�8:V�h�����V�����Q�ec�����N�y�E4���ߺ�x�o��t�����L�F��,#{�BK
 4x�j���������^�,k.��n瞰"o`�}�` ��?�vHc������EM���� R��@/!����Y�� �k�*C����Sچr���b(�@&hx��S#�}��mF�M(d�6������aM�x|{p�B�J�ݱ�/��[�IS��:5J���x���Tl��r]�gf°EY�o4��n�9�aGp�9d+D	n���:w�3�R��]0��Թr*h�HjMO��V6��u��Ԇ0;���?�Ӊ僚	|�˥3
~e�K��Vz�#+Pc���d�IkM^�/jc���o�cPk�������������P�������5�ޣ�|�mu�dg3���7L�Q%�	]�h����d_gw�sM��Mi+�Z�c�/�d=u��"�>��۲��58:F����Y�ﺷ�aε�:+% Z�c<�?�����,��ʎM�p��l�ǈTV7$z��ԯ�J:ᯂ���*���o��˓��.Վ~�t�~����Q~Y��\����YU�*�W�얺�P�q�\�b/C�"�w�L7����E}+ݟ�!���	�)�<p*o%XB��u�Y�P��i�)j:9;�FF�HRo���5�tq��H��cu�z�q�Lĩ��A�Ol��$2��d+=�x��B��S$3�seEtu�,8'��u�$���qL����a�2!�t��O����U�seg _�o�gdv���i
L��-�Q%����`���vi9`g����e�>�ݜ�s�.�n�Ì�wn�n���-U���7����K[�^��q��f��z�?��ꄄP������t��=QHF����a�ZpJdy�ZY��|��RL��ms|�s^O�s��9P;m���G�E��w�#�A��Q�d��7@��[G��ur3 E4���]2|�wo���O�oC�N���*�v��`s����f�:�a��%���ssUOƟ	���F�7�FܰkA#<���Q{m�.o��
'*�8
�fCN�]ia-E7�s���uM�Mm/�.��S���컓R�Vm�G������}u����C$������eO�;��s�/_iH]?������u-���O���-쨕a���s�m�:��5�8��h����TCo�895�˙Hо9��a+}H:���nl#
���Jh`�d'��]�H�t�)�;�B=�3������Xxn����1o�p�����ejת��Y ���.7I"Hʮ J��T&�稝�H{?9�8�c��}@�#��N6�K����E��EC�,���{������5~i��~>t�&K3e���P�p�^s����\��I����?v����Lr6��Y����N�k��/vd�smi�a��t�d��f�U91�c�((h������ �=D2I�%��LvgU��йXV�ֲ"2;Q�n����a��03	�B�亙ƛQu�.4J��)�810ߔ���oK#����Y�ro�iЛ����o	� tY'�W��\�����I� �A��G��𝥞\,�5�zO*�����\&Ȉt^�G�pg�b�	��_#xȺ��dZ\}O�9�"��B��K�?L$/���L�τM�13ż<�������oSP<�/��N:�㠻��<�S��޷�i�j��{K�o��@�S�{�k�)ڰQ�m�+����y���,wD�1o/^itd��|��N$�3���Mp=���{|��(��2,�uc4IY	��*��dSl���3r����6�y��mKGIh�̟|����-2�L\h�n{��ҟ;���lֱ16�.4��уj,R=�"�{a~�h��/�X*�®���B�N$~މ�*Ϝk�<��?�'4g�K,�,��9f;I�@J,�}�Z�7�ݹ�&�L�Ӭe���G�G0�d^�	l�aUec���s���H�y ��j��H��I�<��%g�����˽�|2�����rO��������2[�#�BjL�d�wO��3����"gȋ"�������[��\?���e�FFn��-�vd�jW��ZIf�jeJv��ш>c��D {���cķ-�I���OQ�>T^4Խt�g$�6�" +;w�q�X��Y�l�W�Qq<�Zd� tpA�[@�k�"�O�2whE1�ׇ������Շ�ˀ��e�T�����,*YU�H�|C �}��d������RLYX��؍�4�C���9^<,bԉq��/��f&��\�.�O�ޚ#��TL����j9㣿�Q���a#VM�����I�k��k� ]<ZRD�dqF T-0>J�2f)���z��?�'E7yj�a���.�M��ϣ���B4vT0*M��':.�qy{گ�
Ɗ����W�1o۴����W��򫖝���/�v���)�&�ʈFY=���z�$�.�"�0�{ě����1�*���į���<t�J��!���t<�'�v�3f&՘�칗�'�ɒ�ZGO���:�_ i�뿳~A-�:�ǟ~��9�Llm�eAɶƕh�W��gz$��V3��Xz MQMmi�8��E�9b��$9��ʿ������c�;	���td�
��(�Ҧ��6�m��dò�T�j��I�XIW=Up;^��T� J��x-[PD�,�E�iHy�#e��~^�� -B崥�ǝ�֓v�M�,2�	z@-_3�mB��H��@3xڸ�����]wE��-�2D�	�CH C�3��U��܎@���u2�����,�"x]�u?77��Z�{ðЩ��C�9� �-р
���%����#Htj9��c\������^���Ycd���Z���� YH�\�������ք^�	��%(�W>`\�5���ܸ��^�1z`�I����R�ps�xl~r��xʌ��|#�T�I�hs_0�&�l��GP�	�o!B�K�0OiG���fD��ۮx^w^CF^{�`���i��|�-mfX��i�a�?��s�Fzw*�MU?`f�%��~��g���c<�t;XR�Z@���BZW�`.����S��#��j��輩Q���⼁D��#Ti�S�qڤ?9B�/)���q�*F�-�Q.k��o���q��͡�*q�7#���-'Px Hq�CeG^�1�oA��d�^��ۣ�(Ѿ�}��#�V�
�1���u��^�(���<�;�����JM��S���>�&�V��&�Q)�Ǒ�V �Aj�ŉL�ZW��x�]��������\�d0Z�j�z=��ǿcc)�ڸ�Ø|�֛$5~��z�,���'q�?ўZ�a���!�,�^�܁�6Z_�Z��Ie,<:^�����?pR���x7{�vǌ�;�Eu�,#,�j��X�<*Q� �ǎ�Xs68ϋœ���Z��7Iu�/����JQi�e�3E.b�{�A\F�wo��9���c�`vq\F.GG�;���3�������iLN�av�f��#�!jv�hNa�Q�Y��z�d�ڄR'��`�s�}B��R��30U]1v��:pA}T<�<sO�f���{l@@Q6wU�C'����QJ�:���,�Z ���>��zo@2`�A��,g�=a�>O�V�<������Z����uP���L���g)�?��7y�4w5z0��q|�U���&=�~h�����ыو��i�a[ז�@���-��H��=�C<6e,�����f�
�_#+r������W�K �i!tq�e�X�����/ ��ٜ����x=�<��{EQ�f$JKz�ε��\Hp <=��c�'SKp�C�>El��ԝnl�O�ؖ=D��*���r.A����������^44������@��L�X��BB�^y�]u��	��u����	ѵ�8����ܖ@�~�L0�T3�T�&�P���It�k���/m8LM���R��U����=Rg�&���6�<Ϫp0�w~S
h��C<:�<¢�F ��Q�@�H.v^�$�����%�1S���w������o�
"5�o%���z�/��=�y���ۚ�oa�'1$� �1�B��a��ZQh��$��F�;�9�QNf�2]�����Y�ѳ�ƥ��q���#u�UD	�9m�Y�t�������˲P*�hC��[�\&�c��R�c��%������:�/���q�����;�a�����G��8�	��y��/�}�p��-����t�O>�������j���N�
z2��ӻ'2y8I�@���:���v��C{K=L�����bw�F?(gl�xgd����X�;v����X:�C�����Ȳ#ge*7@`Pd <�kg��f�N�˕�ڪ$��E�*� Bm`2���w2����­F��\ȢAME7 �}����	]�G�n�.���˚���[%��h��^R����4k��	S)���9l��=h�%�A$�Q� ^���J���-hC��Mq�,���R=�!�6�jf�TeJ��o�Ά�G�OF��N}�.�3�.�U[�S1��!���jK+�v���i�;\�mI���\"d��,UY��B1Q��{��4�<^A�������G�Ǒ���\bn���JP�x�)���E"G�r��ZJ7��R��9���\ ���u��7�A�@��:��gD��G�����!�Ve�i61�q{��*xt�C|�ph�nY�~���7#-�a�T��&�n���w�Q�,�_*?2��6���P<�Sǲy}p���y,c �d��%�y��Hl ��tL��;w��$�`*v�j���ExU�0J�/��e{���m�G��"�S��4.�1�9\>��Čl?��'&���D��#�_���%Dg��|Ak�����eiҿ�I�G��oa������}���vz�st0�Eg���^kT[�Jr�8 ����S��_Ag�0�;;��k��u�Px��N	����h���ъ��+�`��u���x'x��e�r�ʶ]�n��㲠AF �
;�Cge	�:�]D�IR[�K���O=�'3��и���A�D�RXP��8�-,�*���'��A�k ?�����\��?��@U�<o1��)p�����#�"D^�)����ǆ,�,y�E?��)�����(]^gu�5R�|�#�#k*D��|�� j��*3����t�M<h�t���S�����X)�R�A�}e4յn�%Ƥ��`1˥�bhDD�{����L�=�X�c]�:�@�Cc��/�b���i�1���ѝ8>o�R�Rأ�&y�� $�*4�Z��˙t�1���ÿyC�r�*�k��$���GRc������� 奇���1b����?��~��|�<�����hv�a���:��A��3{`yZ����3n�ΐy��y|�����k��/e/���F3�n6�/�`R�aP1���B���G!����9��]�0LC����p��}#Z�I"��ylQv���̶��j�yљ�>�����xp��)��-�/��\I����8)r���oJļv N� fy�j�l(TSA��
�g�ޞ����|L��4�E#�ś��p���$�l#P�m'W��N�s`@��@�(i����Q��P]��r��0aWT�;��ݝ	���U+�$�ֲV9���g��l����ᙩ�l>w���2�4����2���Z ��_ng��{jn}�w<}	L%[G0l���Ob_أ���e�]j��'F�"�(2�~�l2le�sRe��kH�X�%;fPzuѕ�PT߆��H
E�_D��� ����	���9��{�?�h�L	�)��R�r��De;5�����L�����y"<�{+ rY-iY��Wg�\!�&@���W�� x��df�Ԩ��(�O=����Չ/&�ߘ�M�i����(#o!��	!/�����;��f��1��bcym-���������@f��f�j:�:�n2�_�J�ޗ����r�wC�g�Y�����Y��ʀ	թ�.5�9�p#��ŷ�&��ms��o��I�/���A�UoU)�;����x�.@wsYN���]c��0������XY�9�m�R��W�A0Jf2��G0(d����w7�R~ǜ�D)�d��v�(�Sd����EnsT�xtPfX�J$�'����WQ��O�!N�?v�m
�����SІT�v���=�A�5_R��e{A� �S�z�� ��QR=.�
>)��(��*5:"�!�!�l|W� ��/+D�Kq)˛�P7V�KFl%��X�YjZ��N��W	jR��X��){y$$��=���&D��\/e=�H���GM
5C�����(f�����O@f��[iK�󥸸�yV ��w��)&�*hE��Ƭ?���IS�1����a݋[�����F�b3�G�Uß�95���e]��Ռ͔ƣE��.�
�\I)r�������x-Ҵ�h��rv�Z9sx�.Qns�%q%����l魫�T1����������� h`gw�Q�Ew��$��?v������Pp�,��(G�)�����W
��k9 w���9Yo|�F%L=s�<`����4\J�����`��b�!����MD>�{��.ǻf��AD������'�d���K��� {,�� ��^=���J��g_�jG�M�����m�@��{�Ĭk�;�ϳ#�>�����ҏ��eЏ9��&ukC?���cD}�����zo&,ty����yP_�qca���g�X�h������o�|��)����0��k�&�:q�NjGl�Q.J�!��گ�&O�.y�3�����F;�L.% �o��Z���Ƹ�N�+OrL!9A�΢�P�cch�GR�i6�~ǥ�������4�
R��	��T�u^��h�#޻[X?���S�F�;p��ȍ���]O9YUk��A����=��I)Z�������;�P���^A��;�B��z,�y,�g�*��`��B6r�ϩ��#�1q�v�燓��t����%\���������4f���8,0��&�&k�N�OB1X���#ߌ��0B���A�����g��b��!?gW"�xyq6������E����(���g�9�����w�8��g���A�Y���^!H!q10"\�m��P��K�Z��,��&f\�#
��yZ�y� ��L��;�A䚪,�������N:6,�P�iF�x
i����(X/x4J|����dv�U`O��uq�_����H0n�O��S����b@P_�V-�`�9d	��-&୪�!���"���e��B>�0C�^Z3g��� ���dI�I���݊z�C*J��o*_�q7�B�e �2{���؞�"+>�wH��+�_?����6�)���`W�R�5�mR�R�~�k���P�)>0bV�ȗ	���.H��h�[8 ��=:�0ad��}��� ���bE�z6s��m���c�[�3Њ�{Ů�f'b��eٝ,���ͼ��}&�X�Â���UeAZ����K/��o�n�iA%�F=�)����*M�!'�S~�+��i<d��%>���Jui
j��yĩ����r�'+�[��ob�Zl�@D�;�W�b u��E���j��ͪ2�F�!6\����UN ��a�*�~H�R���u�˺Bt�N��CL��
���n�XG�P��=wÍ�ϛ.��n�I'4Uw3PMJ
��n���-7ץCE�>rTP�)���5��1���}�c;�nׄ�7w�lR�U�[l���]s?��c��iT��AH�5�����;֚�c";;�~��7��hM�f�Fa��3Wy\^����CYי~��x�L����8RC��1RTM�f����B=O3�8l�B���
Tg-e������R,�.`ƀ������&��^��b�k�ߏR�e���(=��g.�\��X�@�K��s��SGhj�`͑��y����SDJ�cτ�Ͱ�|}��e�ł��
�b���V��)�����
�oȕN�1��-����\�â��Z.��͊-�$�$IC_郟�KX4����:�D�M�����(���JP�ρ8Q���b�C>I��1ز���ЀZ�o�|?���ņ�<�m薎����*�d�Q�����=�}L_'#��U.\�կ��(��.B���a��l�	VT�ݐ�u��f��,�D��k�����Jg���K�su��#��{YN1�R���[T��K�\Y��!n�H(�U��3Lߞ��!C�q:����3"����@?��ء%ޱ���[WN�k�U�)�º!�O=�6���F��p����$s�0�~ 0���yW>�w?�8t��e�jji�7��*��t��3��G�2?|wxCd,�=��,'px��)�r�/J��h�3�@���^C���jE��EԸ��.0��lT���>�N�0(aW�nw����HΑ�zV����*V����N�>8S�����Gޫ�6���)�>�^���C *�āS[�3$0l���|Pg�}쫬����7k��v�m����O\z@1Χ��(#)��#�����-�������Zo��(�����+B�>R�L%��g`�S���I�ږ���^��I^n��;�rM_We���%B�0P1q��'�?=2���ک�W^��$�!<w�/�ݍf�x�� �����.��ѝ]���A�� ���R�t?���Y��=�r�;FF���j?���g!\�?�C[����96e-���ePp��s;z��xNB����2�b��:ǆr@���֏��X\��ݤ��1�t)Ua�< e4 ��E9f���?�g��Z���+��[agŋ�ر��{]��F����"$Fڿ�q��
���͊Az�HnT�z����oTX�-��%�:r�*�$���_%!c�A'i�Az9�Ѫ#&B&,	U4� l�hl|�͜oL܃��sꏸ�Q�J�G�{�(�ZB��#A\���r��A���&�g]�Fk8��ˀ��£��f��(4��Q�+�X�/�d�w�S��0��Y��B@��Kb�hE�_����o�F��������6��F��&Ŋ���ň�3t��)�N�ܖ���Wl�eXu'y��q@|I�+���h�'�"�2HM5�D��Jn:F�4߄��"���c�Q�$�ɼ��^��g+8�cbЃc��7: ��O�d��7,�3��q#%Ʃ
��O��-�f��O:�=7:HS��Ng���@#Q�ڎ��ΦI�*sm����+��^�0��w[�=j��n=<)�t9S�h�C�)S�"%� 4#[�2%��G2G d֬`h��]�K7�9�����1 �e�'��$ⓟ���ѳtqRJ��4��`n@X�(^ Y4a;:�e��HEx���7��(�s�xKA!�!\"y�0�PL?3�HVK�����K_�����~��%AJnD�!["+;ɵ�\@�\$XX"�=E�]Qz�#�6�i^^K�K�弘k��3���z��e���䞏�I�2=������\��	�ʡEx����ۥ�� �-��dd��w,�9��sb�Rˈ�x���S��O�"��.���i�~~��<��������r����kZ䙼�!*W����CS�Y'�N���+�SC�xV2RHS@�߆F�����P�胐k��A���2��uBj��Y��1d���]��V����(��#����elr������bv0D�������
q�c������И�[:�����=��,��������f:vk����̩Q$<�jj�)h��y�L�Xg��6�(�D兂vJ[��G>Jم7d�݅55�3�S�[v�������|JШ]�x�[�r
k����H���,)ߵ#�-�wO��G|<���.}H�4� ?fx�A�H�8�<�1/7`�ɂY�X�:d�����2��b�k���cM;T����A��I���-44E��v'O�5ͭ|B�0�i���|W��9�g
 �䅅�G��]G� �5�rX'�$�8�όa.��m�g��O䶞	��ܔ~y����'<�������_*���T��N�dp������ �ѵd31R'�CjCAL_. >?"2K�E*�8}�Iu@����0V���7���4v��9?�L����Á_%a��}"�?ND	@�Z?+GL?�X�x�kp�|�uӴ�[Q���p�r!��OKLN�-�?�݌5�|��3�FBDB��׏F���&l�F�ե3�����%�y������ۖ���R�rQT�z�lzkT�G���|���@��;��E1�Q&��$,��j�D�*�s̎^*�f�L����;m�3`��$H)�*O���Ka�U$�>�Vk�jE�V��m�Re>��F/�ئ��
������f!Lޤ�3��L��-�;Zs��6	z�1*�Ừ�	Q\jm�β��V�����ʠX�w����/�d�������m�ρx[������?��k !�7���YX�IQ����.4�������6A�Ċ����� �,�c%?)���0M���o>�M1�<�b�?�4�<S>� �({,צ{\�C�M�:,R�N��� 	����^�Z��ۋ��]"�q��d���o:�F�y�u6�;08<C*k
�ayeIR0r6`�M�Nx����8:U���芅hO��)�#lBF�V�������48ض��`Mƭ��e��ڞm|�1�~�2k.���@c.�`�p�ȜC4��=�KX�Ï�8<�J�i��2-'�����d��0g�v�o�Y��,�U��*�LO>�wο����D��>��c���4�]u0,��"�^��qcT?W�rv�W�;b�v��`˶X S��������?�q�D4"H{�$�	���4?�0?�m���m�#s���b��.0�Pω G�BG��*]�ߛU�@?�M�
Wx�'t�B`$]���ק��.�%1�����/-W�/+���AГƯ2 |��Lg�)�
��ݧe
oџ���M볕�Ί�ZK4�)�����Az ϴZ��ĳE��!o��D�@)晟��c���OIL������Y���b��K�h:����Ck-	{�I��)l0XT�eA�H���N&�	�k�M��M��[%(�tR����n�����	`��,d8�^�g?ٕd�o�rϏ�(ؿ(�I��L'Y��	��\�}��xE����.w����9��UMd���`9￀0A�Ar�I�8�s�G���n�UČ$�yM���^c0������}��V<�p����vw�uE`1U�j#Y�z�&�bT��e�t)���d���k�`K�qc�H<�ν���=4��x�F��>��/l4�l�,!��r]���ju<$���%bË:��CO}��&���ΙZ��"�&�	�^��C�XP�雴�՘p��Jd�X��º�}7C�f���d��@RL7���.�ˤ$[S�E.+�SԞI�QO�[�d�qQ�ט�K9��Hg�Di� ����)+
��J���G(�!+oGQ6�>� ��F�v�77�pO�l���r�֣ �oo"W7�h� =Z�d�XAV�g<��O9��x���X/�U�-�v{qJ���*D=}��q�vqa�ۄ����hf�N��מY����?)�i�I��}�Tm(�?�l<�W����DO����-@��n����F�A}%���{����[-!_�p�4�{��#�ƶ�#��1MR�Xh�@}��.&+ �a8��>�P���L�N�*Op�g��R�� ��1O���ߟ��^
q���K�(r̼ʉ�3е�rN���8݀��5�b��W4�å��M~筁����/�I��ʃ��16��
DjP�,�FދO%h�A��}��ڜ��l�`�/m������v{��/BB�>*�'�*<�f��� D�ِB���&`$�uo���Mu�����/H���p$-�G�����a���A�x��~ù���/�F�8�,ݶ�LM��Y:�A?0E�
�+qY�
�ךv`^g��ג7�
����)���l,������u�n	���#C5���y�d���Ҁ�B���I�&)���A;�ny(���Z%S�7�n�#+I��8Z׮��L�9T9�`�Z��3�3���*�k]4"��	�%$3ɠ�G^c/g��b���#�� 8�b���S�As|���n���?��GH��ׯ?&�{�����i�c�x�^^�^Kt#pgF��("t�v��i(�b��	���E��
����Y���r��K"Pze5�r��;������LQ�2�̷.q0����>�>��*9D!�m �'噾A�.G_��1$ge���8�v�,��(n�c���l����&퐗��ɧ ��f&����wg@I�A٤�, �ځ�=�Po/�UBϓ�҉�P'�$%i�|gz�촿�S�ntf�%ܩP��9G��!�µp7`��͒?�S��N��`*f}�h���	�p|o���0�xٌC�8D ��r��n��_,�݉�=��F�T��b4��]a��W��0�U��u������]�eP8ے���o�̀���!\�>����I��%q�I�^.b�!-��܈�my"\m�Sfl	�w��p|�A�A�#o�wc�j&�4���B��3:|�~5��}4����p�%AyT7�7Y��"��r`�H�s�N�j@���Cm�����@��O��@^q �w��)޻���c
>f�X�ڿVw-1����4�ɑM����e:V|/�,g��tW�	6����;6� i	�V�zq��O�}�v^:0+A`[̲t_�汉��7�̂����Jsos،�B���rMF�!F���nW�b�}���m����25�z���i!�++Q���t=�,"qp�	ɏ��^j��0s�&�s�g*�a���8�qW7�߹E���_����Qw����RRP7��<N��d"�ٌ��{�X���Kv��%���-A��b�Ϟ9`2j,:�r���$*�X#q���4�A��IN��Y'{�4�7f:c�!�)����\����Q0<��Ԝ ��N,��Y�Z�sR-`s�rk2F�]��o$��H��ۭGA:2a�o+���0��Ȗ�~ov�r��!Pl[���
�Q��n�[j�g���G]��(=�������8�-R�d>m�kZNmu�/�ru�tS�Y��j�9R���Ziժ�/ag��FJ�C�M������y Ŵ������XFn�[�d䧾�4*CS*	�TC�����9�D���qz���f0C�c�B���Y�wl��)M`����1	�zj�r^[+�#w�M�+C��ނGd��-��:^��䦂;"y����~��GʙY7���u�Wt�|/��:\$������|�.����$��K+�]'B�=�J�:�5{��"�z�J{X#%A6ALQ0ݵv����ߣy�2�����4�@�(���{~.[݃�(��4����/�G�˳
r�B�� ��2V�2�.TK}F���t�D[����u�!�<�ڽ6np��K$U5]�N�Е �>GlZ8{��l�T��~��J���3�)�Q��� ���2Qj�8h��zv��0r ���`��2�l;n�aM*�d�9��S��<*�Ѡ>!J��}rz�G�h˅�w�|3a/�i2�e��j��_��h��}��Qi��0�	ȝ�a;����'��-��'!^�ߑ�J�q�f1F���}��$]�qӝ�B@sW�Mq����3&TK��ynx5B�z��ґi����p<�!���$�nf[�<LHP#��WB�$�_n3��H�R�o�HR#���jE�9���wl�4���E�������I�6o+���>���S젳�qQ�	�qߐ��46(�����ϼ�r9L�V��^�1�r�d�ܖ\�k�s^Ƨ� &
�5R}G���P�s4��LUA��D'r(py_��J�*�u��-�o褐PH)D�(&�����x=��˾;=��5�roc�����E0���.mBx�q
B�!���Ƥc����_,��m7'���P�@׶���������5���+-�隘@F2�w���#��=&����+���R�k�ZѴi��Ϗ�?�u����nv�4�T(�k�$3�K��ЊW��i��� �5E�\�g���N�ܰ1v���*��-*`Z�	���~�,Ùy�i�EU�>A�S��g>;D�vPմ������%��s�%�;>�5���m�ܜnF�sz��{:�H�)��8�ܫ��O��+��;�\�(c4�&����w��:G�N������8b�g=i�z�~m�(�W���5l��� l]M}��O�r
�>s:%<x���#�}[t�yW��qjj:����s/�:Nԯ�B�qjF�Լ$�� �<T�� �z�Id�L�Yyْ$~�a�����}Ï�#o�e�BR�|��G
��Y0܆����V�IѢ��p�qrN��(��4L��<�Cp��h� �u��K�Sp���7��e�^�1��y�+Hsn���K7x9M�{O��	�<DƝE� 2-��mM`Wܷ��	0*�x��h��~���*'��JK�P1 ������{��k��kiP����#��!�
�j��z��nt*�qM���"/��al,�&�ɍ��2E�|��}Vf����{�����m�Ōȏ�ȵ>Y� �u~��Z\p�-�(��X�0<�#�V_��]L	O �9��9=�
'�(�]Ȕ_��ڂ���]�K,���Z�(��M���&��ޙ�%��뽽�W�ڡq� Jj����4��b*�K���v���D����=J�D��'m���2�^]����>&F����B�6%_g������ﳜt-�N���^jd�,��b$���P����f�n�U�+w�W�����14���5F-:d�/�;�d��f��_8�1r��uY��1����B�+���@ز~5�΍#Bl}$%E�T�Ջ��Q�Й��k>���RO�R��U��qC��Z$����t4�B)K]4l��S��qM�}�i	�	\��E"}��<v���·���SA���@��Π�ٟd�@Hz�����3��4�l�W�K�?U�s�\4�|3R�G����JdyOE�����_�����y�ژ��7Doq��L݄D���e��"����W�F�ej��s�z�DRT!�y����Uj03��E�X�I kS���棤�u�F���g�9���(�7��|�:=6�����^���7�)����g��{c����	�u�-������>;���/�-�a@O���-�-m��o���XPYʲ� ��Q���^8��ώ��	6^�1؏�`�H��4A�T���rY���|���7�`���{������}{�5p���`�c�>�1Y�Zy^�Y�X�Y����d.�,�/�p�r���Gk+*����B��ݵ|O�4��$^:߰���p�����2~TKb��Fo:2�"���O�)A�0�)W��k�UO��T�&rW f��]�<��g�E{o�e�8����#�)q�p�~u	��R$Rg:2sb�|�k�@�p�F���\5�V�A/���:[�L�����	��7V��F�DEMHҋa5nϻ�Jt�`s�fq�t��U:sr��6b�F�}P���?�{҆�զ��k��)$1� ��J�{�?��Q8B��'�Mx%YӈI�����N&� 0%�	i]ZwX���`ǗNXM�����55�۷zA�j����u�jt�Ȑ�^v�<��_x)!�~�}5��K��Zr'Hz������KǂǠji�X<���E�@VgY����`"(`�+�<v�;����e��q�o ��޹\��-I��q�Bj���吒v��r�*�8B�]c�oN�2�������p0o�=Thk��X2d�G�q�L�'F��!g=�����SOA�H���h����$����
�ю��cI�r�ևn����2��ߠ�_@��s0}ʁ^8V���aH�	%�v���敽?t��|`��S5��.��/8�A�z5D�^ReE��$�Dǭ\����:HI������Wҝ��3���#���~?(����l����A.�6�}ó�����r	��x�F45x"��V�Η�`�h���2����T2�-������G�u�m9��G�����F@�Saj�	�i��w�ڶ_T��P���d:���k�B�E@��P����@s���e}����z�e,�%6Mo\�]n� �`
(��2�\^Hx�C2�t�
�y��e��Ġ��x��(��Qp~5�N'uR4�鴹�I�uԿ��Ѓſ0q��ԟ�W5�d?�2�¿�&W~��G��c��Hc_	�5���qfP�@R����@KR��.i�Qx�ÕSf���ξ�jG6�;8�P�@y���fV���f��Cp������c��i��&M$�P�Y&��_{�C���sOp��-Qҷ�`���a!ϋ ��U�l����,W/>? Q~��Ӣ��,1��&�k�p�%�{.N�mt�7{Y�,�O��@�$,�A}�d�Mc��'�IYO3|W��$�������{�V��	��Cޯ���WG��d_�� *�5���'Կ�y��E��D�쐾ct" ��M�����خ����'�*��DS�Ϯ"w,��H�{�=���Vi���W��i+|�ɺ�Gs�^Fw�lx��"x�Rn��ìK4�M����Xri�#r�o?L`J�t���5���n��l�5�%x�.��荛�>{�
���Γ�1Ljw�EV���O^���L���_*̚�t�>���׬D�U�p��M�kZ��e5��NT��ǌU��x������eni�7�b�jl���
B�!�9����!8��v@y ����]��F��/�e
{S��U�3�s\�#�q���]���s�C]!�:ܿ#l�G',R�O��}��e��l%%�ކ��B�R�|��?'���B= !��Η�2��3��P�J�h��#������Pm��H�6F��W�.������EO��O����3~:<�eXE^�FT���dj��� ��[<gD����ʐ�`�u��`E��YM��6�%����0��q�ҳ��<T�Q���I��������p���v��n��� ���MC�݀R���#��> (NC!}���\b��J��/��?L
T��E�0"�a_�I=�1�j��C�)6�#B��J�A��aj�W
�¨�Xb�3�;��r�I�|� �~�v�6�4Ķ%u�>�f8 ;��	x�HV~���y� A�O�1��t�nT>osD �|�ƹ*�C}��.�Y��oNd�N�t��V;�^�%%�+��%�d�/j�»ί���}�X�n?�b� ؼ`�X�3'������e�AV��ui܇�E�}X���>c�e��4P@��B�J_����.S���rI�d]�b��{�*��ƍ �B��Xߙ�]���H:���v@_+�u�m�M�k��\�6E��T�ims�9wI���&Ӊ�
�گ��ͭTrG�*�pV�$E��,���(�8�ܲ{$|�ĝ�����8�A���]	��gwt|�F��m̅ Z6����0Z�C�B���ρ8�By���l�Ѭ�FX2���b�~k�'Ì�tS1�[���ϵn,��2����!�CuTO�E�#��x����1���hfYwLKpV�]@���7j�J�ڭ?k	$z��_� ���̝+Q_Eċ��t�ݛl]�]�_���)�<#�FJ����v�3HM��N�ƒռ��J��g�,ڥH���7��ee�*O���i#��-E�p��?�r���=�E�����wd%��z��@��Qk���jt��Ң��;�jx�֑�v}f0.���Y��q���&?&�?I��أ�jp
��!�p��7%�	@��ڹ�jc�ޑsH�Sc	�Y��Y��-<]�U<�R;A��:H����C�!u#��m-݊�R��%�`��jZ����^ e-}�����U�p�N�)UV�Tft�Jv���-Y
�3�A�}n�)��ot �k�..4� �I�-$EAU���ͭ���@�M�D���u�/E�*�7�H^ܣQ� ܠ�+aM<MA�wj	���'�_x�DS�N��>�7o��A��1�xb���=6��ꍃ���mh��z�V�+\���'������r��yL��%cTj����$���닧KD��D�cP�!�6��0QJ���Qg!��f�ߑ��NW�eۊЖ�^���~��#��pG���P���:���Ľv��8���y�A��[����z�R���׸����/in�4(]�a�����kBGS�@��ԸX�{���D00��'�b.�{:}F�$���,�]\3��x�Uŋ鰮oVs7,�_��)^w*\*uk�ʼ��$�����;�ٓT�Q�U��E�?d��5���bB!C>�4�N���,��:�-��M\W�H5��U)Q��ۓG����6Z�w�Dp���������"�Fוd�ܺ��4�u�/*�Wd���`�v��ƚ�R�*�e����(v ����*�}Mi}F��| x0~���Q#�;�|�dt��\W����O�0�����[�̀���7�'�i�X��er%Q�mԥ��r<*(��o�ȧ2�" �[�[�ư}m�(6���c�}���$�#*�d��h��u܃�}�n3ks�_b#��f���VMu3rQ�s�����-Q�%�]��a*H����;5�m��V�6*e lc�6���'0��0v)��6�mW��7�:�i�����5`V[�/-���o(� `�A�HH�l��y0�����9̀��g@}21dO@h4�Eo4�Iaa��b�N��� �ɦ�Z(JA���( ����:%c�Mr�Iی�P�}���,9�dx�aQ��|����`�d1�^;�o�~N4�j���[9[���S�rɻG��{����Äݵ>�c �'2���^�67b;�J�1ʵX�!Y��8�I1�K����T�1G�ϥ�=F����1+{�N�FO���(�Ϲ���}$�q9|���ޤo�F��LI�H���j݊a[(���M=�~nUR��Ջ�ݲ`Ù���y�A�����bH�"Ԩʜ!��'t��{yW�w���@]9�Cn3�F7&ܱv����(�8�g���d�.�JzN#��]�N6�:��n��e���	{��2�~1C�")�8��2����%���/�Q�{!?���J�V�mg�lX�S>A���t}P����H.-6K݃������R�l�/�D����t�3Lk���8^J�s��ą��k���Bj��rýJ���+&l��؊y�dβ
DArǿz��W(_ӈ���.��0���S� 6%�=������bcX�����8SU�t��O|d���mř	h)B$.�7ÅӈGj�%�I�]����!�Pc����X�����7?�1��"1��0��x��3�Ӂ�f��"A���&�z|��bn�R��񔛉�8�R
��������$ �n&�i��̕�N�_�J���z��40/#y����
��1��_��Bnrkf��s�S��b�����K�xX� v�d�W�2wEcG�U:���?��O}��ރ��qd�DK�0o�1�P?<  ��I�:��W�_{h��C���V�QY*^q�:�<��t������6�7�|���!�P��*�}D���|�u;��&��Q��N:����d쳫���hF�<aj'���HKjY�٠t-�,�1&|o�zT�HagB��y���zH�@�O�ͧ�C����LN�_$j�u�+xF߁���p��Xq��u�89.�md�P��"�:�ҬR-h���%i�S_�4K\5\����d-��:e��ɩ�?�%�P���C�.�F�z7�9���A��e7�,c��f4A�6��rE7�l�;�0�e��r�̎��:��=.=``=R#|4��s��O�Z����C��,�F�`~*�
 ���|���01�<n�M���L�aQ��`�˫U�k�_ThH\�B��6�[+����g�(n��F`=v�z�Tɍ�&�ɞt��b�e:�1!��#A��i�ojԂ֦���K�ï��rN_�ȉ�`������Fp�5�Sn[x��|�P�hT�r���=~?�H����f6��pu��֪�	���:2E��7�D����U�TG0|+ن��~?�VC�*��k��&�I㫎�)o��Sx��LkBp����.C����-�){��B ���)S<�]���A�p%,=�پ�����#ф�f��4e8��k!��A�m��������A�ի{�A�K����?�n	Q.�UW�*�ΕN)M�o�`���A�,n2p'{&�����k�M�L��T��!�e��>@�Ac�p���� �����Д
���I��]WR�/{WEg�E���=���_j����\g�5�[}7�[��,��̡w+��
p����p��'��%bĐ7���]{f��I�,? 3�J
VK���t�$b
�2 �w�:$��"��l�Q���
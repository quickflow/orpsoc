// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II"
// VERSION "Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Full Version"

// DATE "11/03/2009 12:35:42"

// 
// Device: Altera EP3C5F256C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module altera_ddr (
	local_address,
	local_write_req,
	local_read_req,
	local_burstbegin,
	local_wdata,
	local_be,
	local_size,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n,
	local_ready,
	local_rdata,
	local_rdata_valid,
	reset_request_n,
	mem_cs_n,
	mem_cke,
	mem_addr,
	mem_ba,
	mem_ras_n,
	mem_cas_n,
	mem_we_n,
	mem_dm,
	local_refresh_ack,
	local_wdata_req,
	local_init_done,
	reset_phy_clk_n,
	phy_clk,
	aux_full_rate_clk,
	aux_half_rate_clk,
	mem_clk,
	mem_clk_n,
	mem_dq,
	mem_dqs)/* synthesis synthesis_greybox=1 */;
input 	[22:0] local_address;
input 	local_write_req;
input 	local_read_req;
input 	local_burstbegin;
input 	[31:0] local_wdata;
input 	[3:0] local_be;
input 	[1:0] local_size;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;
output 	local_ready;
output 	[31:0] local_rdata;
output 	local_rdata_valid;
output 	reset_request_n;
output 	[0:0] mem_cs_n;
output 	[0:0] mem_cke;
output 	[12:0] mem_addr;
output 	[1:0] mem_ba;
output 	mem_ras_n;
output 	mem_cas_n;
output 	mem_we_n;
output 	[1:0] mem_dm;
output 	local_refresh_ack;
output 	local_wdata_req;
output 	local_init_done;
output 	reset_phy_clk_n;
output 	phy_clk;
output 	aux_full_rate_clk;
output 	aux_half_rate_clk;
inout 	[0:0] mem_clk;
inout 	[0:0] mem_clk_n;
inout 	[15:0] mem_dq;
inout 	[1:0] mem_dqs;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[2] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[3] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[4] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[5] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[6] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[7] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[8] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[9] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[10] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[11] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[12] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[13] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[14] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[15] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cs_n[0].cs_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cke[0].cke_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[0].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[1].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[2].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[3].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[4].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[5].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[6].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[7].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[8].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[9].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[10].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[11].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[12].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[0].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[1].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ras_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cas_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|we_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|ddio_outa[0]~dataout ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_n|auto_generated|ddio_outa[0]~dataout ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[2] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[3] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[4] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[5] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[6] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[7] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[8] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[9] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[10] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[11] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[12] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[13] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[14] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[15] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[0] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[1] ;
wire \altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ready~combout ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|locked~combout ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|local_refresh_ack~combout ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[0]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[1]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[2]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[3]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[4]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[5]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[6]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[7]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[8]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[9]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[10]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[11]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[12]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[13]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[14]~q ;
wire \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[15]~q ;
wire \~GND~combout ;
wire \mem_clk[0]~input_o ;
wire \mem_clk_n[0]~input_o ;
wire \mem_dqs[0]~input_o ;
wire \mem_dqs[1]~input_o ;
wire \local_read_req~input_o ;
wire \local_write_req~input_o ;
wire \local_burstbegin~input_o ;
wire \global_reset_n~input_o ;
wire \pll_ref_clk~input_o ;
wire \soft_reset_n~input_o ;
wire \local_address[10]~input_o ;
wire \local_address[16]~input_o ;
wire \local_address[22]~input_o ;
wire \local_address[15]~input_o ;
wire \local_address[19]~input_o ;
wire \local_address[8]~input_o ;
wire \local_address[18]~input_o ;
wire \local_address[21]~input_o ;
wire \local_address[11]~input_o ;
wire \local_address[17]~input_o ;
wire \local_address[9]~input_o ;
wire \local_address[14]~input_o ;
wire \local_address[20]~input_o ;
wire \local_address[13]~input_o ;
wire \local_address[12]~input_o ;
wire \local_be[2]~input_o ;
wire \local_be[0]~input_o ;
wire \local_be[3]~input_o ;
wire \local_be[1]~input_o ;
wire \local_size[0]~input_o ;
wire \local_size[1]~input_o ;
wire \local_address[0]~input_o ;
wire \local_address[1]~input_o ;
wire \local_address[2]~input_o ;
wire \local_address[3]~input_o ;
wire \local_address[4]~input_o ;
wire \local_address[5]~input_o ;
wire \local_address[6]~input_o ;
wire \local_address[7]~input_o ;
wire \local_wdata[16]~input_o ;
wire \local_wdata[0]~input_o ;
wire \local_wdata[17]~input_o ;
wire \local_wdata[1]~input_o ;
wire \local_wdata[18]~input_o ;
wire \local_wdata[2]~input_o ;
wire \local_wdata[19]~input_o ;
wire \local_wdata[3]~input_o ;
wire \local_wdata[20]~input_o ;
wire \local_wdata[4]~input_o ;
wire \local_wdata[21]~input_o ;
wire \local_wdata[5]~input_o ;
wire \local_wdata[22]~input_o ;
wire \local_wdata[6]~input_o ;
wire \local_wdata[23]~input_o ;
wire \local_wdata[7]~input_o ;
wire \local_wdata[24]~input_o ;
wire \local_wdata[8]~input_o ;
wire \local_wdata[25]~input_o ;
wire \local_wdata[9]~input_o ;
wire \local_wdata[26]~input_o ;
wire \local_wdata[10]~input_o ;
wire \local_wdata[27]~input_o ;
wire \local_wdata[11]~input_o ;
wire \local_wdata[28]~input_o ;
wire \local_wdata[12]~input_o ;
wire \local_wdata[29]~input_o ;
wire \local_wdata[13]~input_o ;
wire \local_wdata[30]~input_o ;
wire \local_wdata[14]~input_o ;
wire \local_wdata[31]~input_o ;
wire \local_wdata[15]~input_o ;


altera_ddr_altera_ddr_controller_phy altera_ddr_controller_phy_inst(
	.dq_datain_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[0] ),
	.dq_datain_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[1] ),
	.dq_datain_2(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[2] ),
	.dq_datain_3(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[3] ),
	.dq_datain_4(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[4] ),
	.dq_datain_5(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[5] ),
	.dq_datain_6(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[6] ),
	.dq_datain_7(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[7] ),
	.dq_datain_8(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[8] ),
	.dq_datain_9(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[9] ),
	.dq_datain_10(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[10] ),
	.dq_datain_11(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[11] ),
	.dq_datain_12(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[12] ),
	.dq_datain_13(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[13] ),
	.dq_datain_14(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[14] ),
	.dq_datain_15(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[15] ),
	.q_b_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ),
	.q_b_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ),
	.q_b_2(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ),
	.q_b_3(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ),
	.q_b_4(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ),
	.q_b_5(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ),
	.q_b_6(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ),
	.q_b_7(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ),
	.q_b_16(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ),
	.q_b_17(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ),
	.q_b_18(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ),
	.q_b_19(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ),
	.q_b_20(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ),
	.q_b_21(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ),
	.q_b_22(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ),
	.q_b_23(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ),
	.q_b_8(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ),
	.q_b_9(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ),
	.q_b_10(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ),
	.q_b_11(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ),
	.q_b_12(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ),
	.q_b_13(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ),
	.q_b_14(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ),
	.q_b_15(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ),
	.q_b_24(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ),
	.q_b_25(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ),
	.q_b_26(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ),
	.q_b_27(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ),
	.q_b_28(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ),
	.q_b_29(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ),
	.q_b_30(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ),
	.q_b_31(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ),
	.clk_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[0] ),
	.clk_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[1] ),
	.dataout_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cs_n[0].cs_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_01(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cke[0].cke_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_02(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[0].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_03(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[1].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_04(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[2].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_05(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[3].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_06(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[4].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_07(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[5].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_08(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[6].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_09(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[7].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_010(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[8].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_011(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[9].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_012(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[10].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_013(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[11].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_014(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[12].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_015(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[0].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_016(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[1].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_017(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ras_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_018(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cas_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_019(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|we_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ),
	.dm_ddio_dataout_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[0] ),
	.dm_ddio_dataout_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[1] ),
	.ddio_outa_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|ddio_outa[0]~dataout ),
	.ddio_outa_01(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_n|auto_generated|ddio_outa[0]~dataout ),
	.dq_ddio_dataout_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[0] ),
	.dq_ddio_dataout_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[1] ),
	.dq_ddio_dataout_2(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[2] ),
	.dq_ddio_dataout_3(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[3] ),
	.dq_ddio_dataout_4(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[4] ),
	.dq_ddio_dataout_5(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[5] ),
	.dq_ddio_dataout_6(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[6] ),
	.dq_ddio_dataout_7(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[7] ),
	.dq_ddio_dataout_8(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[8] ),
	.dq_ddio_dataout_9(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[9] ),
	.dq_ddio_dataout_10(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[10] ),
	.dq_ddio_dataout_11(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[11] ),
	.dq_ddio_dataout_12(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[12] ),
	.dq_ddio_dataout_13(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[13] ),
	.dq_ddio_dataout_14(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[14] ),
	.dq_ddio_dataout_15(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[15] ),
	.dqs_ddio_dataout_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[0] ),
	.wdp_wdqs_oe_2x_r_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[0] ),
	.dqs_ddio_dataout_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[1] ),
	.wdp_wdqs_oe_2x_r_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[1] ),
	.ready(\altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ready~combout ),
	.ctl_rdata_valid_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ),
	.reset_request_n(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|locked~combout ),
	.ctl_init_success(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ),
	.local_refresh_ack(\altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|local_refresh_ack~combout ),
	.reset_phy_clk_1x_n(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ),
	.wdp_wdata_oe_2x_r_0(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[0]~q ),
	.wdp_wdata_oe_2x_r_1(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[1]~q ),
	.wdp_wdata_oe_2x_r_2(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[2]~q ),
	.wdp_wdata_oe_2x_r_3(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[3]~q ),
	.wdp_wdata_oe_2x_r_4(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[4]~q ),
	.wdp_wdata_oe_2x_r_5(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[5]~q ),
	.wdp_wdata_oe_2x_r_6(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[6]~q ),
	.wdp_wdata_oe_2x_r_7(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[7]~q ),
	.wdp_wdata_oe_2x_r_8(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[8]~q ),
	.wdp_wdata_oe_2x_r_9(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[9]~q ),
	.wdp_wdata_oe_2x_r_10(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[10]~q ),
	.wdp_wdata_oe_2x_r_11(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[11]~q ),
	.wdp_wdata_oe_2x_r_12(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[12]~q ),
	.wdp_wdata_oe_2x_r_13(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[13]~q ),
	.wdp_wdata_oe_2x_r_14(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[14]~q ),
	.wdp_wdata_oe_2x_r_15(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[15]~q ),
	.GND_port(\~GND~combout ),
	.mem_clk_0(\mem_clk[0]~input_o ),
	.local_read_req(\local_read_req~input_o ),
	.local_write_req(\local_write_req~input_o ),
	.local_burstbegin(\local_burstbegin~input_o ),
	.global_reset_n(\global_reset_n~input_o ),
	.pll_ref_clk(\pll_ref_clk~input_o ),
	.soft_reset_n(\soft_reset_n~input_o ),
	.local_address_10(\local_address[10]~input_o ),
	.local_address_16(\local_address[16]~input_o ),
	.local_address_22(\local_address[22]~input_o ),
	.local_address_15(\local_address[15]~input_o ),
	.local_address_19(\local_address[19]~input_o ),
	.local_address_8(\local_address[8]~input_o ),
	.local_address_18(\local_address[18]~input_o ),
	.local_address_21(\local_address[21]~input_o ),
	.local_address_11(\local_address[11]~input_o ),
	.local_address_17(\local_address[17]~input_o ),
	.local_address_9(\local_address[9]~input_o ),
	.local_address_14(\local_address[14]~input_o ),
	.local_address_20(\local_address[20]~input_o ),
	.local_address_13(\local_address[13]~input_o ),
	.local_address_12(\local_address[12]~input_o ),
	.local_be_2(\local_be[2]~input_o ),
	.local_be_0(\local_be[0]~input_o ),
	.local_be_3(\local_be[3]~input_o ),
	.local_be_1(\local_be[1]~input_o ),
	.local_size_0(\local_size[0]~input_o ),
	.local_size_1(\local_size[1]~input_o ),
	.local_address_0(\local_address[0]~input_o ),
	.local_address_1(\local_address[1]~input_o ),
	.local_address_2(\local_address[2]~input_o ),
	.local_address_3(\local_address[3]~input_o ),
	.local_address_4(\local_address[4]~input_o ),
	.local_address_5(\local_address[5]~input_o ),
	.local_address_6(\local_address[6]~input_o ),
	.local_address_7(\local_address[7]~input_o ),
	.local_wdata_16(\local_wdata[16]~input_o ),
	.local_wdata_0(\local_wdata[0]~input_o ),
	.local_wdata_17(\local_wdata[17]~input_o ),
	.local_wdata_1(\local_wdata[1]~input_o ),
	.local_wdata_18(\local_wdata[18]~input_o ),
	.local_wdata_2(\local_wdata[2]~input_o ),
	.local_wdata_19(\local_wdata[19]~input_o ),
	.local_wdata_3(\local_wdata[3]~input_o ),
	.local_wdata_20(\local_wdata[20]~input_o ),
	.local_wdata_4(\local_wdata[4]~input_o ),
	.local_wdata_21(\local_wdata[21]~input_o ),
	.local_wdata_5(\local_wdata[5]~input_o ),
	.local_wdata_22(\local_wdata[22]~input_o ),
	.local_wdata_6(\local_wdata[6]~input_o ),
	.local_wdata_23(\local_wdata[23]~input_o ),
	.local_wdata_7(\local_wdata[7]~input_o ),
	.local_wdata_24(\local_wdata[24]~input_o ),
	.local_wdata_8(\local_wdata[8]~input_o ),
	.local_wdata_25(\local_wdata[25]~input_o ),
	.local_wdata_9(\local_wdata[9]~input_o ),
	.local_wdata_26(\local_wdata[26]~input_o ),
	.local_wdata_10(\local_wdata[10]~input_o ),
	.local_wdata_27(\local_wdata[27]~input_o ),
	.local_wdata_11(\local_wdata[11]~input_o ),
	.local_wdata_28(\local_wdata[28]~input_o ),
	.local_wdata_12(\local_wdata[12]~input_o ),
	.local_wdata_29(\local_wdata[29]~input_o ),
	.local_wdata_13(\local_wdata[13]~input_o ),
	.local_wdata_30(\local_wdata[30]~input_o ),
	.local_wdata_14(\local_wdata[14]~input_o ),
	.local_wdata_31(\local_wdata[31]~input_o ),
	.local_wdata_15(\local_wdata[15]~input_o ));

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[0]  = mem_dq[0];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[1]  = mem_dq[1];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[2]  = mem_dq[2];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[3]  = mem_dq[3];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[4]  = mem_dq[4];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[5]  = mem_dq[5];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[6]  = mem_dq[6];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[7]  = mem_dq[7];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[8]  = mem_dq[8];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[9]  = mem_dq[9];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[10]  = mem_dq[10];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[11]  = mem_dq[11];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[12]  = mem_dq[12];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[13]  = mem_dq[13];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[14]  = mem_dq[14];

assign \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_datain[15]  = mem_dq[15];

cycloneiii_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

assign \mem_clk[0]~input_o  = mem_clk[0];

assign \local_read_req~input_o  = local_read_req;

assign \local_write_req~input_o  = local_write_req;

assign \local_burstbegin~input_o  = local_burstbegin;

assign \global_reset_n~input_o  = global_reset_n;

assign \pll_ref_clk~input_o  = pll_ref_clk;

assign \soft_reset_n~input_o  = soft_reset_n;

assign \local_address[10]~input_o  = local_address[10];

assign \local_address[16]~input_o  = local_address[16];

assign \local_address[22]~input_o  = local_address[22];

assign \local_address[15]~input_o  = local_address[15];

assign \local_address[19]~input_o  = local_address[19];

assign \local_address[8]~input_o  = local_address[8];

assign \local_address[18]~input_o  = local_address[18];

assign \local_address[21]~input_o  = local_address[21];

assign \local_address[11]~input_o  = local_address[11];

assign \local_address[17]~input_o  = local_address[17];

assign \local_address[9]~input_o  = local_address[9];

assign \local_address[14]~input_o  = local_address[14];

assign \local_address[20]~input_o  = local_address[20];

assign \local_address[13]~input_o  = local_address[13];

assign \local_address[12]~input_o  = local_address[12];

assign \local_be[2]~input_o  = local_be[2];

assign \local_be[0]~input_o  = local_be[0];

assign \local_be[3]~input_o  = local_be[3];

assign \local_be[1]~input_o  = local_be[1];

assign \local_size[0]~input_o  = local_size[0];

assign \local_size[1]~input_o  = local_size[1];

assign \local_address[0]~input_o  = local_address[0];

assign \local_address[1]~input_o  = local_address[1];

assign \local_address[2]~input_o  = local_address[2];

assign \local_address[3]~input_o  = local_address[3];

assign \local_address[4]~input_o  = local_address[4];

assign \local_address[5]~input_o  = local_address[5];

assign \local_address[6]~input_o  = local_address[6];

assign \local_address[7]~input_o  = local_address[7];

assign \local_wdata[16]~input_o  = local_wdata[16];

assign \local_wdata[0]~input_o  = local_wdata[0];

assign \local_wdata[17]~input_o  = local_wdata[17];

assign \local_wdata[1]~input_o  = local_wdata[1];

assign \local_wdata[18]~input_o  = local_wdata[18];

assign \local_wdata[2]~input_o  = local_wdata[2];

assign \local_wdata[19]~input_o  = local_wdata[19];

assign \local_wdata[3]~input_o  = local_wdata[3];

assign \local_wdata[20]~input_o  = local_wdata[20];

assign \local_wdata[4]~input_o  = local_wdata[4];

assign \local_wdata[21]~input_o  = local_wdata[21];

assign \local_wdata[5]~input_o  = local_wdata[5];

assign \local_wdata[22]~input_o  = local_wdata[22];

assign \local_wdata[6]~input_o  = local_wdata[6];

assign \local_wdata[23]~input_o  = local_wdata[23];

assign \local_wdata[7]~input_o  = local_wdata[7];

assign \local_wdata[24]~input_o  = local_wdata[24];

assign \local_wdata[8]~input_o  = local_wdata[8];

assign \local_wdata[25]~input_o  = local_wdata[25];

assign \local_wdata[9]~input_o  = local_wdata[9];

assign \local_wdata[26]~input_o  = local_wdata[26];

assign \local_wdata[10]~input_o  = local_wdata[10];

assign \local_wdata[27]~input_o  = local_wdata[27];

assign \local_wdata[11]~input_o  = local_wdata[11];

assign \local_wdata[28]~input_o  = local_wdata[28];

assign \local_wdata[12]~input_o  = local_wdata[12];

assign \local_wdata[29]~input_o  = local_wdata[29];

assign \local_wdata[13]~input_o  = local_wdata[13];

assign \local_wdata[30]~input_o  = local_wdata[30];

assign \local_wdata[14]~input_o  = local_wdata[14];

assign \local_wdata[31]~input_o  = local_wdata[31];

assign \local_wdata[15]~input_o  = local_wdata[15];

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[0].dm_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[0] ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[0]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[0].dm_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[0].dm_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[1].dm_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm_ddio_dataout[1] ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[1]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[1].dm_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dm[1].dm_obuf .open_drain_output = "false";

assign local_ready = \altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ready~combout ;

assign local_rdata[0] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ;

assign local_rdata[1] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ;

assign local_rdata[2] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ;

assign local_rdata[3] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ;

assign local_rdata[4] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ;

assign local_rdata[5] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ;

assign local_rdata[6] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ;

assign local_rdata[7] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ;

assign local_rdata[8] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ;

assign local_rdata[9] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ;

assign local_rdata[10] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ;

assign local_rdata[11] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ;

assign local_rdata[12] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ;

assign local_rdata[13] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ;

assign local_rdata[14] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ;

assign local_rdata[15] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ;

assign local_rdata[16] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ;

assign local_rdata[17] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ;

assign local_rdata[18] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ;

assign local_rdata[19] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ;

assign local_rdata[20] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ;

assign local_rdata[21] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ;

assign local_rdata[22] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ;

assign local_rdata[23] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ;

assign local_rdata[24] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ;

assign local_rdata[25] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ;

assign local_rdata[26] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ;

assign local_rdata[27] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ;

assign local_rdata[28] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ;

assign local_rdata[29] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ;

assign local_rdata[30] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ;

assign local_rdata[31] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdp|full_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ;

assign local_rdata_valid = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ;

assign reset_request_n = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|locked~combout ;

assign mem_cs_n[0] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cs_n[0].cs_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_cke[0] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cke[0].cke_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[0] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[0].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[1] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[1].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[2] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[2].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[3] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[3].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[4] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[4].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[5] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[5].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[6] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[6].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[7] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[7].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[8] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[8].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[9] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[9].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[10] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[10].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[11] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[11].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[12] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|addr[12].addr_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ba[0] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[0].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ba[1] = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ba[1].ba_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ras_n = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|ras_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_cas_n = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|cas_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_we_n = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|full_rate_adc_gen.adc|we_n_struct|full_rate.addr_pin|auto_generated|dataout[0] ;

assign local_refresh_ack = \altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|local_refresh_ack~combout ;

assign local_wdata_req = gnd;

assign local_init_done = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ;

assign reset_phy_clk_n = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ;

assign phy_clk = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[1] ;

assign aux_full_rate_clk = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[1] ;

assign aux_half_rate_clk = \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|pll|altpll_component|auto_generated|clk[0] ;

cycloneiii_io_obuf \mem_clk[0]~output (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|ddio_outa[0]~dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_clk[0]),
	.obar());
defparam \mem_clk[0]~output .bus_hold = "false";
defparam \mem_clk[0]~output .open_drain_output = "false";

cycloneiii_io_obuf \mem_clk_n[0]~output (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].ddr_clk_out_n|auto_generated|ddio_outa[0]~dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_clk_n[0]),
	.obar());
defparam \mem_clk_n[0]~output .bus_hold = "false";
defparam \mem_clk_n[0]~output .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[0] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[0]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[0]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[1] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[1]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[1]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[2] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[2]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[2]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[3] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[3]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[3]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[4] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[4]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[4]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[5] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[5]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[5]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[6] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[6]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[6]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[7] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[7]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[7]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[8] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[8]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[8]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[9] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[9]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[9]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[10] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[10]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[10]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[11] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[11]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[11]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[12] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[12]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[12]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[13] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[13]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[13]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[14] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[14]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[14]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dq_ddio_dataout[15] ),
	.oe(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdata_oe_2x_r[15]~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[15]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[0].dqs_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[0] ),
	.oe(!\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[0] ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[0]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[0].dqs_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[0].dqs_obuf .open_drain_output = "false";

cycloneiii_io_obuf \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[1].dqs_obuf (
	.i(\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs_ddio_dataout[1] ),
	.oe(!\altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|wdp_wdqs_oe_2x_r[1] ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[1]),
	.obar());
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[1].dqs_obuf .bus_hold = "false";
defparam \altera_ddr_controller_phy_inst|altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|dpio|dqs[1].dqs_obuf .open_drain_output = "false";

assign \mem_clk_n[0]~input_o  = mem_clk_n[0];

assign \mem_dqs[0]~input_o  = mem_dqs[0];

assign \mem_dqs[1]~input_o  = mem_dqs[1];

endmodule

module altera_ddr_altera_ddr_controller_phy (
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dm_ddio_dataout_0,
	dm_ddio_dataout_1,
	ddio_outa_0,
	ddio_outa_01,
	dq_ddio_dataout_0,
	dq_ddio_dataout_1,
	dq_ddio_dataout_2,
	dq_ddio_dataout_3,
	dq_ddio_dataout_4,
	dq_ddio_dataout_5,
	dq_ddio_dataout_6,
	dq_ddio_dataout_7,
	dq_ddio_dataout_8,
	dq_ddio_dataout_9,
	dq_ddio_dataout_10,
	dq_ddio_dataout_11,
	dq_ddio_dataout_12,
	dq_ddio_dataout_13,
	dq_ddio_dataout_14,
	dq_ddio_dataout_15,
	dqs_ddio_dataout_0,
	wdp_wdqs_oe_2x_r_0,
	dqs_ddio_dataout_1,
	wdp_wdqs_oe_2x_r_1,
	ready,
	ctl_rdata_valid_0,
	reset_request_n,
	ctl_init_success,
	local_refresh_ack,
	reset_phy_clk_1x_n,
	wdp_wdata_oe_2x_r_0,
	wdp_wdata_oe_2x_r_1,
	wdp_wdata_oe_2x_r_2,
	wdp_wdata_oe_2x_r_3,
	wdp_wdata_oe_2x_r_4,
	wdp_wdata_oe_2x_r_5,
	wdp_wdata_oe_2x_r_6,
	wdp_wdata_oe_2x_r_7,
	wdp_wdata_oe_2x_r_8,
	wdp_wdata_oe_2x_r_9,
	wdp_wdata_oe_2x_r_10,
	wdp_wdata_oe_2x_r_11,
	wdp_wdata_oe_2x_r_12,
	wdp_wdata_oe_2x_r_13,
	wdp_wdata_oe_2x_r_14,
	wdp_wdata_oe_2x_r_15,
	GND_port,
	mem_clk_0,
	local_read_req,
	local_write_req,
	local_burstbegin,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n,
	local_address_10,
	local_address_16,
	local_address_22,
	local_address_15,
	local_address_19,
	local_address_8,
	local_address_18,
	local_address_21,
	local_address_11,
	local_address_17,
	local_address_9,
	local_address_14,
	local_address_20,
	local_address_13,
	local_address_12,
	local_be_2,
	local_be_0,
	local_be_3,
	local_be_1,
	local_size_0,
	local_size_1,
	local_address_0,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_6,
	local_address_7,
	local_wdata_16,
	local_wdata_0,
	local_wdata_17,
	local_wdata_1,
	local_wdata_18,
	local_wdata_2,
	local_wdata_19,
	local_wdata_3,
	local_wdata_20,
	local_wdata_4,
	local_wdata_21,
	local_wdata_5,
	local_wdata_22,
	local_wdata_6,
	local_wdata_23,
	local_wdata_7,
	local_wdata_24,
	local_wdata_8,
	local_wdata_25,
	local_wdata_9,
	local_wdata_26,
	local_wdata_10,
	local_wdata_27,
	local_wdata_11,
	local_wdata_28,
	local_wdata_12,
	local_wdata_29,
	local_wdata_13,
	local_wdata_30,
	local_wdata_14,
	local_wdata_31,
	local_wdata_15)/* synthesis synthesis_greybox=1 */;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dm_ddio_dataout_0;
output 	dm_ddio_dataout_1;
output 	ddio_outa_0;
output 	ddio_outa_01;
output 	dq_ddio_dataout_0;
output 	dq_ddio_dataout_1;
output 	dq_ddio_dataout_2;
output 	dq_ddio_dataout_3;
output 	dq_ddio_dataout_4;
output 	dq_ddio_dataout_5;
output 	dq_ddio_dataout_6;
output 	dq_ddio_dataout_7;
output 	dq_ddio_dataout_8;
output 	dq_ddio_dataout_9;
output 	dq_ddio_dataout_10;
output 	dq_ddio_dataout_11;
output 	dq_ddio_dataout_12;
output 	dq_ddio_dataout_13;
output 	dq_ddio_dataout_14;
output 	dq_ddio_dataout_15;
output 	dqs_ddio_dataout_0;
output 	wdp_wdqs_oe_2x_r_0;
output 	dqs_ddio_dataout_1;
output 	wdp_wdqs_oe_2x_r_1;
output 	ready;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	ctl_init_success;
output 	local_refresh_ack;
output 	reset_phy_clk_1x_n;
output 	wdp_wdata_oe_2x_r_0;
output 	wdp_wdata_oe_2x_r_1;
output 	wdp_wdata_oe_2x_r_2;
output 	wdp_wdata_oe_2x_r_3;
output 	wdp_wdata_oe_2x_r_4;
output 	wdp_wdata_oe_2x_r_5;
output 	wdp_wdata_oe_2x_r_6;
output 	wdp_wdata_oe_2x_r_7;
output 	wdp_wdata_oe_2x_r_8;
output 	wdp_wdata_oe_2x_r_9;
output 	wdp_wdata_oe_2x_r_10;
output 	wdp_wdata_oe_2x_r_11;
output 	wdp_wdata_oe_2x_r_12;
output 	wdp_wdata_oe_2x_r_13;
output 	wdp_wdata_oe_2x_r_14;
output 	wdp_wdata_oe_2x_r_15;
input 	GND_port;
input 	mem_clk_0;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;
input 	local_address_10;
input 	local_address_16;
input 	local_address_22;
input 	local_address_15;
input 	local_address_19;
input 	local_address_8;
input 	local_address_18;
input 	local_address_21;
input 	local_address_11;
input 	local_address_17;
input 	local_address_9;
input 	local_address_14;
input 	local_address_20;
input 	local_address_13;
input 	local_address_12;
input 	local_be_2;
input 	local_be_0;
input 	local_be_3;
input 	local_be_1;
input 	local_size_0;
input 	local_size_1;
input 	local_address_0;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_6;
input 	local_address_7;
input 	local_wdata_16;
input 	local_wdata_0;
input 	local_wdata_17;
input 	local_wdata_1;
input 	local_wdata_18;
input 	local_wdata_2;
input 	local_wdata_19;
input 	local_wdata_3;
input 	local_wdata_20;
input 	local_wdata_4;
input 	local_wdata_21;
input 	local_wdata_5;
input 	local_wdata_22;
input 	local_wdata_6;
input 	local_wdata_23;
input 	local_wdata_7;
input 	local_wdata_24;
input 	local_wdata_8;
input 	local_wdata_25;
input 	local_wdata_9;
input 	local_wdata_26;
input 	local_wdata_10;
input 	local_wdata_27;
input 	local_wdata_11;
input 	local_wdata_28;
input 	local_wdata_12;
input 	local_wdata_29;
input 	local_wdata_13;
input 	local_wdata_30;
input 	local_wdata_14;
input 	local_wdata_31;
input 	local_wdata_15;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[34] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[32] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[35] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[33] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_rd[0]~combout ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cs_n[0]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[0]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[1]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[2]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[3]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[4]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[5]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[6]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[7]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[8]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[9]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[10]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[11]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[12]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[0]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[1]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ras_n~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cas_n~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|we_n~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_wlat_r[0]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~0_combout ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|Equal6~0_combout ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~1_combout ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~3_combout ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ;
wire \altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_dqs_burst[0]~0_combout ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas4~q ;
wire \altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas3~q ;


altera_ddr_altera_ddr_auk_ddr_hp_controller_wrapper altera_ddr_auk_ddr_hp_controller_wrapper_inst(
	.clk_1(clk_1),
	.q_b_34(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[34] ),
	.q_b_32(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[32] ),
	.q_b_35(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[35] ),
	.q_b_33(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[33] ),
	.q_b_16(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_17(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_18(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_2(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_19(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_3(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_20(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_4(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_21(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_5(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_22(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_6(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_23(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_7(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_24(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_8(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_25(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_9(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_26(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_10(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_27(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_11(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_28(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_12(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_29(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_13(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_30(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_14(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_31(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_15(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.seq_ac_add_1t_ac_lat_internal(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ),
	.ready(ready),
	.ctl_init_success(ctl_init_success),
	.local_refresh_ack(local_refresh_ack),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_rd_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_rd[0]~combout ),
	.cs_n_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cs_n[0]~q ),
	.a_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[0]~q ),
	.a_1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[1]~q ),
	.a_2(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[2]~q ),
	.a_3(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[3]~q ),
	.a_4(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[4]~q ),
	.a_5(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[5]~q ),
	.a_6(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[6]~q ),
	.a_7(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[7]~q ),
	.a_8(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[8]~q ),
	.a_9(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[9]~q ),
	.a_10(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[10]~q ),
	.a_11(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[11]~q ),
	.a_12(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[12]~q ),
	.ba_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[0]~q ),
	.ba_1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[1]~q ),
	.ras_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ras_n~q ),
	.cas_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cas_n~q ),
	.we_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|we_n~q ),
	.control_wlat_r_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_wlat_r[0]~q ),
	.control_doing_wr(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~0_combout ),
	.Equal6(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|Equal6~0_combout ),
	.control_doing_wr1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~1_combout ),
	.control_doing_wr2(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~3_combout ),
	.wd_lat_0(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ),
	.wd_lat_1(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ),
	.wd_lat_4(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ),
	.wd_lat_3(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ),
	.wd_lat_2(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ),
	.control_dqs_burst_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_dqs_burst[0]~0_combout ),
	.dqs_burst_cas4(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas4~q ),
	.dqs_burst_cas3(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas3~q ),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_address_10(local_address_10),
	.local_address_16(local_address_16),
	.local_address_22(local_address_22),
	.local_address_15(local_address_15),
	.local_address_19(local_address_19),
	.local_address_8(local_address_8),
	.local_address_18(local_address_18),
	.local_address_21(local_address_21),
	.local_address_11(local_address_11),
	.local_address_17(local_address_17),
	.local_address_9(local_address_9),
	.local_address_14(local_address_14),
	.local_address_20(local_address_20),
	.local_address_13(local_address_13),
	.local_address_12(local_address_12),
	.local_be_2(local_be_2),
	.local_be_0(local_be_0),
	.local_be_3(local_be_3),
	.local_be_1(local_be_1),
	.local_size_0(local_size_0),
	.local_size_1(local_size_1),
	.local_address_0(local_address_0),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_6(local_address_6),
	.local_address_7(local_address_7),
	.local_wdata_16(local_wdata_16),
	.local_wdata_0(local_wdata_0),
	.local_wdata_17(local_wdata_17),
	.local_wdata_1(local_wdata_1),
	.local_wdata_18(local_wdata_18),
	.local_wdata_2(local_wdata_2),
	.local_wdata_19(local_wdata_19),
	.local_wdata_3(local_wdata_3),
	.local_wdata_20(local_wdata_20),
	.local_wdata_4(local_wdata_4),
	.local_wdata_21(local_wdata_21),
	.local_wdata_5(local_wdata_5),
	.local_wdata_22(local_wdata_22),
	.local_wdata_6(local_wdata_6),
	.local_wdata_23(local_wdata_23),
	.local_wdata_7(local_wdata_7),
	.local_wdata_24(local_wdata_24),
	.local_wdata_8(local_wdata_8),
	.local_wdata_25(local_wdata_25),
	.local_wdata_9(local_wdata_9),
	.local_wdata_26(local_wdata_26),
	.local_wdata_10(local_wdata_10),
	.local_wdata_27(local_wdata_27),
	.local_wdata_11(local_wdata_11),
	.local_wdata_28(local_wdata_28),
	.local_wdata_12(local_wdata_12),
	.local_wdata_29(local_wdata_29),
	.local_wdata_13(local_wdata_13),
	.local_wdata_30(local_wdata_30),
	.local_wdata_14(local_wdata_14),
	.local_wdata_31(local_wdata_31),
	.local_wdata_15(local_wdata_15));

altera_ddr_altera_ddr_phy altera_ddr_phy_inst(
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.dm_ddio_dataout_0(dm_ddio_dataout_0),
	.dm_ddio_dataout_1(dm_ddio_dataout_1),
	.ddio_outa_0(ddio_outa_0),
	.ddio_outa_01(ddio_outa_01),
	.dq_ddio_dataout_0(dq_ddio_dataout_0),
	.dq_ddio_dataout_1(dq_ddio_dataout_1),
	.dq_ddio_dataout_2(dq_ddio_dataout_2),
	.dq_ddio_dataout_3(dq_ddio_dataout_3),
	.dq_ddio_dataout_4(dq_ddio_dataout_4),
	.dq_ddio_dataout_5(dq_ddio_dataout_5),
	.dq_ddio_dataout_6(dq_ddio_dataout_6),
	.dq_ddio_dataout_7(dq_ddio_dataout_7),
	.dq_ddio_dataout_8(dq_ddio_dataout_8),
	.dq_ddio_dataout_9(dq_ddio_dataout_9),
	.dq_ddio_dataout_10(dq_ddio_dataout_10),
	.dq_ddio_dataout_11(dq_ddio_dataout_11),
	.dq_ddio_dataout_12(dq_ddio_dataout_12),
	.dq_ddio_dataout_13(dq_ddio_dataout_13),
	.dq_ddio_dataout_14(dq_ddio_dataout_14),
	.dq_ddio_dataout_15(dq_ddio_dataout_15),
	.dqs_ddio_dataout_0(dqs_ddio_dataout_0),
	.wdp_wdqs_oe_2x_r_0(wdp_wdqs_oe_2x_r_0),
	.dqs_ddio_dataout_1(dqs_ddio_dataout_1),
	.wdp_wdqs_oe_2x_r_1(wdp_wdqs_oe_2x_r_1),
	.q_b_34(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[34] ),
	.q_b_32(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[32] ),
	.q_b_35(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[35] ),
	.q_b_33(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[33] ),
	.q_b_161(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_01(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_171(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_110(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_181(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_210(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_191(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_36(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_201(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_41(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_211(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_51(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_221(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_61(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_231(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_71(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_241(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_81(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_251(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_91(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_261(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_101(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_271(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_111(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_281(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_121(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_291(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_131(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_301(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_141(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_311(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_151(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|g_local_avalon_if:av_if|wfifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.seq_ac_add_1t_ac_lat_internal(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.reset_request_n(reset_request_n),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_rd_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_rd[0]~combout ),
	.cs_n_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cs_n[0]~q ),
	.a_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[0]~q ),
	.a_1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[1]~q ),
	.a_2(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[2]~q ),
	.a_3(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[3]~q ),
	.a_4(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[4]~q ),
	.a_5(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[5]~q ),
	.a_6(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[6]~q ),
	.a_7(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[7]~q ),
	.a_8(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[8]~q ),
	.a_9(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[9]~q ),
	.a_10(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[10]~q ),
	.a_11(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[11]~q ),
	.a_12(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|a[12]~q ),
	.ba_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[0]~q ),
	.ba_1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ba[1]~q ),
	.ras_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|ras_n~q ),
	.cas_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|cas_n~q ),
	.we_n(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|we_n~q ),
	.wdp_wdata_oe_2x_r_0(wdp_wdata_oe_2x_r_0),
	.wdp_wdata_oe_2x_r_1(wdp_wdata_oe_2x_r_1),
	.wdp_wdata_oe_2x_r_2(wdp_wdata_oe_2x_r_2),
	.wdp_wdata_oe_2x_r_3(wdp_wdata_oe_2x_r_3),
	.wdp_wdata_oe_2x_r_4(wdp_wdata_oe_2x_r_4),
	.wdp_wdata_oe_2x_r_5(wdp_wdata_oe_2x_r_5),
	.wdp_wdata_oe_2x_r_6(wdp_wdata_oe_2x_r_6),
	.wdp_wdata_oe_2x_r_7(wdp_wdata_oe_2x_r_7),
	.wdp_wdata_oe_2x_r_8(wdp_wdata_oe_2x_r_8),
	.wdp_wdata_oe_2x_r_9(wdp_wdata_oe_2x_r_9),
	.wdp_wdata_oe_2x_r_10(wdp_wdata_oe_2x_r_10),
	.wdp_wdata_oe_2x_r_11(wdp_wdata_oe_2x_r_11),
	.wdp_wdata_oe_2x_r_12(wdp_wdata_oe_2x_r_12),
	.wdp_wdata_oe_2x_r_13(wdp_wdata_oe_2x_r_13),
	.wdp_wdata_oe_2x_r_14(wdp_wdata_oe_2x_r_14),
	.wdp_wdata_oe_2x_r_15(wdp_wdata_oe_2x_r_15),
	.control_wlat_r_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_wlat_r[0]~q ),
	.control_doing_wr(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~0_combout ),
	.Equal6(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|Equal6~0_combout ),
	.control_doing_wr1(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~1_combout ),
	.control_doing_wr2(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_doing_wr~3_combout ),
	.wd_lat_0(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ),
	.wd_lat_1(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ),
	.wd_lat_4(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ),
	.wd_lat_3(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ),
	.wd_lat_2(\altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ),
	.control_dqs_burst_0(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|control_dqs_burst[0]~0_combout ),
	.dqs_burst_cas4(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas4~q ),
	.dqs_burst_cas3(\altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller_inst|dqs_burst_cas3~q ),
	.GND_port(GND_port),
	.mem_clk_0(mem_clk_0),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

endmodule

module altera_ddr_altera_ddr_auk_ddr_hp_controller_wrapper (
	clk_1,
	q_b_34,
	q_b_32,
	q_b_35,
	q_b_33,
	q_b_16,
	q_b_0,
	q_b_17,
	q_b_1,
	q_b_18,
	q_b_2,
	q_b_19,
	q_b_3,
	q_b_20,
	q_b_4,
	q_b_21,
	q_b_5,
	q_b_22,
	q_b_6,
	q_b_23,
	q_b_7,
	q_b_24,
	q_b_8,
	q_b_25,
	q_b_9,
	q_b_26,
	q_b_10,
	q_b_27,
	q_b_11,
	q_b_28,
	q_b_12,
	q_b_29,
	q_b_13,
	q_b_30,
	q_b_14,
	q_b_31,
	q_b_15,
	seq_ac_add_1t_ac_lat_internal,
	ready,
	ctl_init_success,
	local_refresh_ack,
	reset_phy_clk_1x_n,
	control_doing_rd_0,
	cs_n_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	ba_0,
	ba_1,
	ras_n,
	cas_n,
	we_n,
	control_wlat_r_0,
	control_doing_wr,
	Equal6,
	control_doing_wr1,
	control_doing_wr2,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	control_dqs_burst_0,
	dqs_burst_cas4,
	dqs_burst_cas3,
	local_read_req,
	local_write_req,
	local_burstbegin,
	local_address_10,
	local_address_16,
	local_address_22,
	local_address_15,
	local_address_19,
	local_address_8,
	local_address_18,
	local_address_21,
	local_address_11,
	local_address_17,
	local_address_9,
	local_address_14,
	local_address_20,
	local_address_13,
	local_address_12,
	local_be_2,
	local_be_0,
	local_be_3,
	local_be_1,
	local_size_0,
	local_size_1,
	local_address_0,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_6,
	local_address_7,
	local_wdata_16,
	local_wdata_0,
	local_wdata_17,
	local_wdata_1,
	local_wdata_18,
	local_wdata_2,
	local_wdata_19,
	local_wdata_3,
	local_wdata_20,
	local_wdata_4,
	local_wdata_21,
	local_wdata_5,
	local_wdata_22,
	local_wdata_6,
	local_wdata_23,
	local_wdata_7,
	local_wdata_24,
	local_wdata_8,
	local_wdata_25,
	local_wdata_9,
	local_wdata_26,
	local_wdata_10,
	local_wdata_27,
	local_wdata_11,
	local_wdata_28,
	local_wdata_12,
	local_wdata_29,
	local_wdata_13,
	local_wdata_30,
	local_wdata_14,
	local_wdata_31,
	local_wdata_15)/* synthesis synthesis_greybox=1 */;
input 	clk_1;
output 	q_b_34;
output 	q_b_32;
output 	q_b_35;
output 	q_b_33;
output 	q_b_16;
output 	q_b_0;
output 	q_b_17;
output 	q_b_1;
output 	q_b_18;
output 	q_b_2;
output 	q_b_19;
output 	q_b_3;
output 	q_b_20;
output 	q_b_4;
output 	q_b_21;
output 	q_b_5;
output 	q_b_22;
output 	q_b_6;
output 	q_b_23;
output 	q_b_7;
output 	q_b_24;
output 	q_b_8;
output 	q_b_25;
output 	q_b_9;
output 	q_b_26;
output 	q_b_10;
output 	q_b_27;
output 	q_b_11;
output 	q_b_28;
output 	q_b_12;
output 	q_b_29;
output 	q_b_13;
output 	q_b_30;
output 	q_b_14;
output 	q_b_31;
output 	q_b_15;
input 	seq_ac_add_1t_ac_lat_internal;
output 	ready;
input 	ctl_init_success;
output 	local_refresh_ack;
input 	reset_phy_clk_1x_n;
output 	control_doing_rd_0;
output 	cs_n_0;
output 	a_0;
output 	a_1;
output 	a_2;
output 	a_3;
output 	a_4;
output 	a_5;
output 	a_6;
output 	a_7;
output 	a_8;
output 	a_9;
output 	a_10;
output 	a_11;
output 	a_12;
output 	ba_0;
output 	ba_1;
output 	ras_n;
output 	cas_n;
output 	we_n;
output 	control_wlat_r_0;
output 	control_doing_wr;
output 	Equal6;
output 	control_doing_wr1;
output 	control_doing_wr2;
input 	wd_lat_0;
input 	wd_lat_1;
input 	wd_lat_4;
input 	wd_lat_3;
input 	wd_lat_2;
output 	control_dqs_burst_0;
output 	dqs_burst_cas4;
output 	dqs_burst_cas3;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	local_address_10;
input 	local_address_16;
input 	local_address_22;
input 	local_address_15;
input 	local_address_19;
input 	local_address_8;
input 	local_address_18;
input 	local_address_21;
input 	local_address_11;
input 	local_address_17;
input 	local_address_9;
input 	local_address_14;
input 	local_address_20;
input 	local_address_13;
input 	local_address_12;
input 	local_be_2;
input 	local_be_0;
input 	local_be_3;
input 	local_be_1;
input 	local_size_0;
input 	local_size_1;
input 	local_address_0;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_6;
input 	local_address_7;
input 	local_wdata_16;
input 	local_wdata_0;
input 	local_wdata_17;
input 	local_wdata_1;
input 	local_wdata_18;
input 	local_wdata_2;
input 	local_wdata_19;
input 	local_wdata_3;
input 	local_wdata_20;
input 	local_wdata_4;
input 	local_wdata_21;
input 	local_wdata_5;
input 	local_wdata_22;
input 	local_wdata_6;
input 	local_wdata_23;
input 	local_wdata_7;
input 	local_wdata_24;
input 	local_wdata_8;
input 	local_wdata_25;
input 	local_wdata_9;
input 	local_wdata_26;
input 	local_wdata_10;
input 	local_wdata_27;
input 	local_wdata_11;
input 	local_wdata_28;
input 	local_wdata_12;
input 	local_wdata_29;
input 	local_wdata_13;
input 	local_wdata_30;
input 	local_wdata_14;
input 	local_wdata_31;
input 	local_wdata_15;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_auk_ddr_hp_controller auk_ddr_hp_controller_inst(
	.clk(clk_1),
	.q_b_34(q_b_34),
	.q_b_32(q_b_32),
	.q_b_35(q_b_35),
	.q_b_33(q_b_33),
	.q_b_16(q_b_16),
	.q_b_0(q_b_0),
	.q_b_17(q_b_17),
	.q_b_1(q_b_1),
	.q_b_18(q_b_18),
	.q_b_2(q_b_2),
	.q_b_19(q_b_19),
	.q_b_3(q_b_3),
	.q_b_20(q_b_20),
	.q_b_4(q_b_4),
	.q_b_21(q_b_21),
	.q_b_5(q_b_5),
	.q_b_22(q_b_22),
	.q_b_6(q_b_6),
	.q_b_23(q_b_23),
	.q_b_7(q_b_7),
	.q_b_24(q_b_24),
	.q_b_8(q_b_8),
	.q_b_25(q_b_25),
	.q_b_9(q_b_9),
	.q_b_26(q_b_26),
	.q_b_10(q_b_10),
	.q_b_27(q_b_27),
	.q_b_11(q_b_11),
	.q_b_28(q_b_28),
	.q_b_12(q_b_12),
	.q_b_29(q_b_29),
	.q_b_13(q_b_13),
	.q_b_30(q_b_30),
	.q_b_14(q_b_14),
	.q_b_31(q_b_31),
	.q_b_15(q_b_15),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ready1(ready),
	.ctl_init_success(ctl_init_success),
	.local_refresh_ack1(local_refresh_ack),
	.reset_n(reset_phy_clk_1x_n),
	.control_doing_rd_0(control_doing_rd_0),
	.cs_n_0(cs_n_0),
	.a_0(a_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.ba_0(ba_0),
	.ba_1(ba_1),
	.ras_n1(ras_n),
	.cas_n1(cas_n),
	.we_n1(we_n),
	.control_wlat_r_0(control_wlat_r_0),
	.control_doing_wr(control_doing_wr),
	.Equal6(Equal6),
	.control_doing_wr1(control_doing_wr1),
	.control_doing_wr2(control_doing_wr2),
	.wd_lat_0(wd_lat_0),
	.control_wlat({wd_lat_4,wd_lat_3,gnd,wd_lat_1,gnd}),
	.wd_lat_2(wd_lat_2),
	.control_dqs_burst_0(control_dqs_burst_0),
	.dqs_burst_cas41(dqs_burst_cas4),
	.dqs_burst_cas31(dqs_burst_cas3),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_row_addr({local_address_20,local_address_19,local_address_18,local_address_17,local_address_16,local_address_15,local_address_14,local_address_13,local_address_12,local_address_11,local_address_10,local_address_9,local_address_8}),
	.local_bank_addr({local_address_22,local_address_21}),
	.local_be_2(local_be_2),
	.local_be_0(local_be_0),
	.local_be_3(local_be_3),
	.local_be_1(local_be_1),
	.local_size({local_size_1,local_size_0}),
	.local_col_addr({local_address_7,local_address_6,local_address_5,local_address_4,local_address_3,local_address_2,local_address_1,local_address_0}),
	.local_wdata_16(local_wdata_16),
	.local_wdata_0(local_wdata_0),
	.local_wdata_17(local_wdata_17),
	.local_wdata_1(local_wdata_1),
	.local_wdata_18(local_wdata_18),
	.local_wdata_2(local_wdata_2),
	.local_wdata_19(local_wdata_19),
	.local_wdata_3(local_wdata_3),
	.local_wdata_20(local_wdata_20),
	.local_wdata_4(local_wdata_4),
	.local_wdata_21(local_wdata_21),
	.local_wdata_5(local_wdata_5),
	.local_wdata_22(local_wdata_22),
	.local_wdata_6(local_wdata_6),
	.local_wdata_23(local_wdata_23),
	.local_wdata_7(local_wdata_7),
	.local_wdata_24(local_wdata_24),
	.local_wdata_8(local_wdata_8),
	.local_wdata_25(local_wdata_25),
	.local_wdata_9(local_wdata_9),
	.local_wdata_26(local_wdata_26),
	.local_wdata_10(local_wdata_10),
	.local_wdata_27(local_wdata_27),
	.local_wdata_11(local_wdata_11),
	.local_wdata_28(local_wdata_28),
	.local_wdata_12(local_wdata_12),
	.local_wdata_29(local_wdata_29),
	.local_wdata_13(local_wdata_13),
	.local_wdata_30(local_wdata_30),
	.local_wdata_14(local_wdata_14),
	.local_wdata_31(local_wdata_31),
	.local_wdata_15(local_wdata_15));

endmodule

module altera_ddr_auk_ddr_hp_controller (
	clk,
	q_b_34,
	q_b_32,
	q_b_35,
	q_b_33,
	q_b_16,
	q_b_0,
	q_b_17,
	q_b_1,
	q_b_18,
	q_b_2,
	q_b_19,
	q_b_3,
	q_b_20,
	q_b_4,
	q_b_21,
	q_b_5,
	q_b_22,
	q_b_6,
	q_b_23,
	q_b_7,
	q_b_24,
	q_b_8,
	q_b_25,
	q_b_9,
	q_b_26,
	q_b_10,
	q_b_27,
	q_b_11,
	q_b_28,
	q_b_12,
	q_b_29,
	q_b_13,
	q_b_30,
	q_b_14,
	q_b_31,
	q_b_15,
	seq_ac_add_1t_ac_lat_internal,
	ready1,
	ctl_init_success,
	local_refresh_ack1,
	reset_n,
	control_doing_rd_0,
	cs_n_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	ba_0,
	ba_1,
	ras_n1,
	cas_n1,
	we_n1,
	control_wlat_r_0,
	control_doing_wr,
	Equal6,
	control_doing_wr1,
	control_doing_wr2,
	wd_lat_0,
	control_wlat,
	wd_lat_2,
	control_dqs_burst_0,
	dqs_burst_cas41,
	dqs_burst_cas31,
	local_read_req,
	local_write_req,
	local_burstbegin,
	local_row_addr,
	local_bank_addr,
	local_be_2,
	local_be_0,
	local_be_3,
	local_be_1,
	local_size,
	local_col_addr,
	local_wdata_16,
	local_wdata_0,
	local_wdata_17,
	local_wdata_1,
	local_wdata_18,
	local_wdata_2,
	local_wdata_19,
	local_wdata_3,
	local_wdata_20,
	local_wdata_4,
	local_wdata_21,
	local_wdata_5,
	local_wdata_22,
	local_wdata_6,
	local_wdata_23,
	local_wdata_7,
	local_wdata_24,
	local_wdata_8,
	local_wdata_25,
	local_wdata_9,
	local_wdata_26,
	local_wdata_10,
	local_wdata_27,
	local_wdata_11,
	local_wdata_28,
	local_wdata_12,
	local_wdata_29,
	local_wdata_13,
	local_wdata_30,
	local_wdata_14,
	local_wdata_31,
	local_wdata_15)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	q_b_34;
output 	q_b_32;
output 	q_b_35;
output 	q_b_33;
output 	q_b_16;
output 	q_b_0;
output 	q_b_17;
output 	q_b_1;
output 	q_b_18;
output 	q_b_2;
output 	q_b_19;
output 	q_b_3;
output 	q_b_20;
output 	q_b_4;
output 	q_b_21;
output 	q_b_5;
output 	q_b_22;
output 	q_b_6;
output 	q_b_23;
output 	q_b_7;
output 	q_b_24;
output 	q_b_8;
output 	q_b_25;
output 	q_b_9;
output 	q_b_26;
output 	q_b_10;
output 	q_b_27;
output 	q_b_11;
output 	q_b_28;
output 	q_b_12;
output 	q_b_29;
output 	q_b_13;
output 	q_b_30;
output 	q_b_14;
output 	q_b_31;
output 	q_b_15;
input 	seq_ac_add_1t_ac_lat_internal;
output 	ready1;
input 	ctl_init_success;
output 	local_refresh_ack1;
input 	reset_n;
output 	control_doing_rd_0;
output 	cs_n_0;
output 	a_0;
output 	a_1;
output 	a_2;
output 	a_3;
output 	a_4;
output 	a_5;
output 	a_6;
output 	a_7;
output 	a_8;
output 	a_9;
output 	a_10;
output 	a_11;
output 	a_12;
output 	ba_0;
output 	ba_1;
output 	ras_n1;
output 	cas_n1;
output 	we_n1;
output 	control_wlat_r_0;
output 	control_doing_wr;
output 	Equal6;
output 	control_doing_wr1;
output 	control_doing_wr2;
input 	wd_lat_0;
input 	[4:0] control_wlat;
input 	wd_lat_2;
output 	control_dqs_burst_0;
output 	dqs_burst_cas41;
output 	dqs_burst_cas31;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	[12:0] local_row_addr;
input 	[1:0] local_bank_addr;
input 	local_be_2;
input 	local_be_0;
input 	local_be_3;
input 	local_be_1;
input 	[1:0] local_size;
input 	[7:0] local_col_addr;
input 	local_wdata_16;
input 	local_wdata_0;
input 	local_wdata_17;
input 	local_wdata_1;
input 	local_wdata_18;
input 	local_wdata_2;
input 	local_wdata_19;
input 	local_wdata_3;
input 	local_wdata_20;
input 	local_wdata_4;
input 	local_wdata_21;
input 	local_wdata_5;
input 	local_wdata_22;
input 	local_wdata_6;
input 	local_wdata_23;
input 	local_wdata_7;
input 	local_wdata_24;
input 	local_wdata_8;
input 	local_wdata_25;
input 	local_wdata_9;
input 	local_wdata_26;
input 	local_wdata_10;
input 	local_wdata_27;
input 	local_wdata_11;
input 	local_wdata_28;
input 	local_wdata_12;
input 	local_wdata_29;
input 	local_wdata_13;
input 	local_wdata_30;
input 	local_wdata_14;
input 	local_wdata_31;
input 	local_wdata_15;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \in_buf|my_fifo|pipefull[3]~q ;
wire \rfsh_counter[10]~q ;
wire \rfsh_counter[3]~q ;
wire \rfsh_counter[5]~q ;
wire \rfsh_counter[15]~q ;
wire \rfsh_counter[11]~q ;
wire \rfsh_counter[3]~54_combout ;
wire \rfsh_counter[5]~58_combout ;
wire \rfsh_counter[10]~68_combout ;
wire \rfsh_counter[11]~70_combout ;
wire \rfsh_counter[14]~77 ;
wire \rfsh_counter[15]~78_combout ;
wire \held_burstbegin~q ;
wire \write_req_to_in_buf~0_combout ;
wire \Selector23~2_combout ;
wire \bank_man|Equal8~0_combout ;
wire \held_burstbegin~2_combout ;
wire \in_buf|my_fifo|pipefull[0]~q ;
wire \in_buf|my_fifo|pipe[0][29]~q ;
wire \Selector0~5_combout ;
wire \in_buf|my_fifo|pipe[0][28]~q ;
wire \Selector0~6_combout ;
wire \ba[1]~117_combout ;
wire \in_buf|my_fifo|pipe[0][27]~q ;
wire \Selector0~7_combout ;
wire \Selector0~8_combout ;
wire \Selector0~9_combout ;
wire \write_req_last~q ;
wire \Selector0~13_combout ;
wire \Selector5~3_combout ;
wire \Selector0~14_combout ;
wire \Selector0~15_combout ;
wire \Selector0~16_combout ;
wire \Selector0~20_combout ;
wire \Selector0~24_combout ;
wire \Selector2~6_combout ;
wire \p_main_fsm~160_combout ;
wire \g_timers:2:bank_timer|twr_pipe[2]~q ;
wire \g_timers:3:bank_timer|twr_pipe[2]~q ;
wire \g_timers:1:bank_timer|twr_pipe[2]~q ;
wire \g_timers:0:bank_timer|twr_pipe[2]~q ;
wire \to_this_bank[2]~q ;
wire \g_timers:2:bank_timer|finished_twr~combout ;
wire \to_this_bank[1]~q ;
wire \g_timers:1:bank_timer|finished_twr~combout ;
wire \to_this_bank[0]~q ;
wire \g_timers:0:bank_timer|finished_twr~combout ;
wire \to_this_bank[3]~q ;
wire \g_timers:3:bank_timer|finished_twr~combout ;
wire \state~329_combout ;
wire \state~330_combout ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \Selector4~3_combout ;
wire \state~331_combout ;
wire \Selector50~0_combout ;
wire \doing_pch_all~q ;
wire \in_buf|my_fifo|pipe[0][9]~q ;
wire \in_buf|my_fifo|pipe[0][8]~q ;
wire \bank_man|Mux11~1_combout ;
wire \bank_man|Mux3~1_combout ;
wire \in_buf|my_fifo|pipe[0][19]~q ;
wire \in_buf|my_fifo|pipe[0][11]~q ;
wire \Equal2~0_combout ;
wire \bank_man|Mux8~1_combout ;
wire \in_buf|my_fifo|pipe[0][14]~q ;
wire \bank_man|Mux2~1_combout ;
wire \in_buf|my_fifo|pipe[0][20]~q ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \bank_man|Mux9~1_combout ;
wire \bank_man|Mux4~1_combout ;
wire \in_buf|my_fifo|pipe[0][18]~q ;
wire \in_buf|my_fifo|pipe[0][13]~q ;
wire \bank_man|Mux12~1_combout ;
wire \bank_man|Mux7~1_combout ;
wire \in_buf|my_fifo|pipe[0][15]~q ;
wire \in_buf|my_fifo|pipe[0][10]~q ;
wire \bank_man|Mux5~1_combout ;
wire \bank_man|Mux6~1_combout ;
wire \in_buf|my_fifo|pipe[0][16]~q ;
wire \in_buf|my_fifo|pipe[0][17]~q ;
wire \Equal2~5_combout ;
wire \bank_man|Mux10~1_combout ;
wire \bank_man|Mux1~1_combout ;
wire \in_buf|my_fifo|pipe[0][21]~q ;
wire \in_buf|my_fifo|pipe[0][12]~q ;
wire \bank_man|Mux0~1_combout ;
wire \in_buf|my_fifo|pipe[0][22]~q ;
wire \bank_man|Mux13~1_combout ;
wire \Selector20~3_combout ;
wire \Selector46~4_combout ;
wire \Selector46~5_combout ;
wire \Selector46~6_combout ;
wire \Selector46~7_combout ;
wire \Selector8~3_combout ;
wire \in_buf|my_fifo|pipe[0][24]~q ;
wire \in_buf|my_fifo|pipe[0][25]~q ;
wire \rdata_bcount_le_1~3_combout ;
wire \wdata_burst_count[1]~52_combout ;
wire \wdata_burst_count[1]~55_combout ;
wire \Selector42~2_combout ;
wire \wdata_burst_count[1]~57_combout ;
wire \wdata_burst_count[1]~58_combout ;
wire \wdata_burst_count[1]~59_combout ;
wire \wdata_burst_count[1]~61_combout ;
wire \wdata_burst_count[1]~62_combout ;
wire \wdata_burst_count[1]~64_combout ;
wire \rdata_bcount_eq_1~2_combout ;
wire \Selector11~0_combout ;
wire \rdata_bcount_eq_0~3_combout ;
wire \Selector43~1_combout ;
wire \Selector43~2_combout ;
wire \Selector45~0_combout ;
wire \Selector45~1_combout ;
wire \dqs_toggle_le_2~q ;
wire \Selector43~4_combout ;
wire \Selector44~4_combout ;
wire \Selector44~5_combout ;
wire \Selector44~6_combout ;
wire \Selector44~7_combout ;
wire \Selector44~8_combout ;
wire \Selector44~10_combout ;
wire \Selector12~3_combout ;
wire \Selector12~5_combout ;
wire \Selector53~7_combout ;
wire \cs_n~60_combout ;
wire \Selector17~0_combout ;
wire \Selector17~1_combout ;
wire \Selector17~4_combout ;
wire \Selector17~7_combout ;
wire \a[0]~577_combout ;
wire \ba[1]~125_combout ;
wire \a[0]~578_combout ;
wire \a[0]~579_combout ;
wire \a[0]~580_combout ;
wire \a[0]~581_combout ;
wire \a[5]~593_combout ;
wire \a[5]~601_combout ;
wire \a[5]~602_combout ;
wire \a[5]~603_combout ;
wire \a[5]~604_combout ;
wire \a[5]~608_combout ;
wire \a[5]~611_combout ;
wire \ba[1]~130_combout ;
wire \ba[1]~131_combout ;
wire \ba[1]~132_combout ;
wire \ba[1]~133_combout ;
wire \ba[1]~134_combout ;
wire \ba[1]~135_combout ;
wire \ba[1]~136_combout ;
wire \ba[1]~137_combout ;
wire \ba[1]~138_combout ;
wire \ba[1]~139_combout ;
wire \ba[1]~140_combout ;
wire \ba[1]~142_combout ;
wire \ba[1]~145_combout ;
wire \ba[1]~146_combout ;
wire \ba[1]~147_combout ;
wire \ba[1]~154_combout ;
wire \ba[1]~155_combout ;
wire \ba[1]~158_combout ;
wire \Selector18~2_combout ;
wire \Selector20~6_combout ;
wire \Selector20~7_combout ;
wire \Selector20~8_combout ;
wire \Selector20~9_combout ;
wire \g_timers:1:bank_timer|finished_tras~q ;
wire \g_timers:2:bank_timer|finished_tras~q ;
wire \g_timers:0:bank_timer|finished_tras~q ;
wire \g_timers:3:bank_timer|finished_tras~q ;
wire \bank_addr_this_valid[1]~q ;
wire \bank_addr_this_valid[0]~q ;
wire \Decoder1~0_combout ;
wire \Decoder1~1_combout ;
wire \Decoder1~2_combout ;
wire \Decoder1~3_combout ;
wire \Selector20~18_combout ;
wire \Selector42~4_combout ;
wire \Selector42~10_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \LessThan0~3_combout ;
wire \LessThan0~4_combout ;
wire \wdata_burst_count[0]~70_combout ;
wire \dqs_toggle_le_2~1_combout ;
wire \in_buf|my_fifo|pipe[0][0]~q ;
wire \in_buf|my_fifo|pipe[0][1]~q ;
wire \in_buf|my_fifo|pipe[0][2]~q ;
wire \in_buf|my_fifo|pipe[0][3]~q ;
wire \in_buf|my_fifo|pipe[0][4]~q ;
wire \in_buf|my_fifo|pipe[0][5]~q ;
wire \in_buf|my_fifo|pipe[0][6]~q ;
wire \in_buf|my_fifo|pipe[0][7]~q ;
wire \Selector0~27_combout ;
wire \Selector42~11_combout ;
wire \Selector46~15_combout ;
wire \Selector12~9_combout ;
wire \ba[1]~162_combout ;
wire \Selector19~9_combout ;
wire \read_req_next~0_combout ;
wire \rfsh_counter[0]~48_combout ;
wire \rfsh_counter[0]~q ;
wire \rfsh_counter[0]~49 ;
wire \rfsh_counter[1]~51 ;
wire \rfsh_counter[2]~53 ;
wire \rfsh_counter[3]~55 ;
wire \rfsh_counter[4]~56_combout ;
wire \rfsh_counter[4]~q ;
wire \rfsh_counter[2]~52_combout ;
wire \rfsh_counter[2]~q ;
wire \rfsh_counter[1]~50_combout ;
wire \rfsh_counter[1]~q ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \rfsh_counter[4]~57 ;
wire \rfsh_counter[5]~59 ;
wire \rfsh_counter[6]~61 ;
wire \rfsh_counter[7]~63 ;
wire \rfsh_counter[8]~65 ;
wire \rfsh_counter[9]~66_combout ;
wire \rfsh_counter[9]~q ;
wire \rfsh_counter[6]~60_combout ;
wire \rfsh_counter[6]~q ;
wire \rfsh_counter[7]~62_combout ;
wire \rfsh_counter[7]~q ;
wire \rfsh_counter[8]~64_combout ;
wire \rfsh_counter[8]~q ;
wire \LessThan1~2_combout ;
wire \LessThan1~3_combout ;
wire \rfsh_counter[9]~67 ;
wire \rfsh_counter[10]~69 ;
wire \rfsh_counter[11]~71 ;
wire \rfsh_counter[12]~72_combout ;
wire \rfsh_counter[12]~q ;
wire \LessThan1~4_combout ;
wire \rfsh_counter[12]~73 ;
wire \rfsh_counter[13]~74_combout ;
wire \rfsh_counter[13]~q ;
wire \rfsh_counter[13]~75 ;
wire \rfsh_counter[14]~76_combout ;
wire \rfsh_counter[14]~q ;
wire \LessThan1~5_combout ;
wire \rfsh_pending~2_combout ;
wire \rfsh_pending~q ;
wire \size_next[1]~1_combout ;
wire \size_this[1]~q ;
wire \accepted_r~q ;
wire \size_last[1]~q ;
wire \Selector37~2_combout ;
wire \bank_is_open~q ;
wire \size_next[0]~0_combout ;
wire \size_this[0]~q ;
wire \size_last[0]~q ;
wire \rdata_burst_count~6_combout ;
wire \rdata_burst_count[0]~q ;
wire \rdata_burst_count~4_combout ;
wire \rdata_burst_count~5_combout ;
wire \rdata_burst_count[1]~q ;
wire \rdata_bcount_eq_1~3_combout ;
wire \rdata_bcount_eq_1~q ;
wire \write_req_next~0_combout ;
wire \write_req_this~q ;
wire \am_writing~25_combout ;
wire \rdata_valid_pipe[3]~q ;
wire \am_reading~0_combout ;
wire \am_reading~q ;
wire \am_reading_r~q ;
wire \Selector50~5_combout ;
wire \p_main_fsm~105_combout ;
wire \Selector5~8_combout ;
wire \state.s_activate~q ;
wire \wdata_burst_count[1]~53_combout ;
wire \wdata_burst_count[1]~54_combout ;
wire \row_addr_next[8]~3_combout ;
wire \row_addr_next[3]~4_combout ;
wire \Equal2~3_combout ;
wire \row_addr_next[5]~5_combout ;
wire \row_addr_next[0]~6_combout ;
wire \Equal2~4_combout ;
wire \row_addr_next[11]~9_combout ;
wire \row_addr_next[2]~10_combout ;
wire \Equal2~6_combout ;
wire \row_addr_next[12]~11_combout ;
wire \Equal2~7_combout ;
wire \Equal2~8_combout ;
wire \this_row_is_open~q ;
wire \wdata_burst_count[1]~63_combout ;
wire \p_main_fsm~19_combout ;
wire \Selector8~2_combout ;
wire \Selector19~6_combout ;
wire \Selector8~4_combout ;
wire \state.s_write~q ;
wire \p_main_fsm~154_combout ;
wire \wdata_burst_count[1]~56_combout ;
wire \wdata_burst_count[1]~51_combout ;
wire \wdata_burst_count[1]~65_combout ;
wire \ba[1]~122_combout ;
wire \wdata_burst_count[1]~60_combout ;
wire \wdata_burst_count[1]~66_combout ;
wire \wdata_burst_count[0]~71_combout ;
wire \wdata_burst_count[0]~q ;
wire \wdata_burst_count[1]~67_combout ;
wire \wdata_burst_count[1]~q ;
wire \rdata_bcount_eq_0~4_combout ;
wire \rdata_bcount_eq_0~q ;
wire \doing_wr_cl_pipe[0]~q ;
wire \finished_twtr~0_combout ;
wire \finished_twtr~q ;
wire \p_main_fsm~158_combout ;
wire \dqs_must_keep_toggling[2]~8_combout ;
wire \dqs_must_keep_toggling[2]~q ;
wire \dqs_must_keep_toggling[0]~7_combout ;
wire \dqs_must_keep_toggling[0]~q ;
wire \dqs_must_keep_toggling[1]~6_combout ;
wire \dqs_must_keep_toggling[1]~q ;
wire \dqs_toggle_le_1~1_combout ;
wire \dqs_toggle_le_1~q ;
wire \Selector20~2_combout ;
wire \rdata_bcount_le_1~4_combout ;
wire \rdata_bcount_le_1~q ;
wire \a[5]~574_combout ;
wire \p_main_fsm~166_combout ;
wire \Selector11~3_combout ;
wire \p_main_fsm~39_combout ;
wire \Selector44~15_combout ;
wire \Selector44~9_combout ;
wire \p_main_fsm~156_combout ;
wire \Selector44~11_combout ;
wire \p_main_fsm~63_combout ;
wire \Selector44~12_combout ;
wire \Selector44~13_combout ;
wire \Selector37~6_combout ;
wire \ba[1]~124_combout ;
wire \Selector37~4_combout ;
wire \Selector37~5_combout ;
wire \didnt_term~q ;
wire \Selector0~28_combout ;
wire \read_req_last~3_combout ;
wire \read_req_last~2_combout ;
wire \read_req_last~q ;
wire \Selector45~2_combout ;
wire \Selector45~3_combout ;
wire \p_main_fsm~61_combout ;
wire \Selector45~4_combout ;
wire \Selector45~5_combout ;
wire \Selector45~6_combout ;
wire \cs_addr_to_term[0]~q ;
wire \ba[1]~121_combout ;
wire \Selector44~14_combout ;
wire \didnt_read~q ;
wire \ba[1]~118_combout ;
wire \Selector43~3_combout ;
wire \Selector43~0_combout ;
wire \Selector10~0_combout ;
wire \row_mux_sel_next[0]~1_combout ;
wire \bank_addr_this[0]~q ;
wire \row_mux_sel_next[1]~0_combout ;
wire \row_mux_sel_last[1]~2_combout ;
wire \buf_not_empty_r~q ;
wire \row_mux_sel_last[1]~3_combout ;
wire \row_mux_sel_last[0]~q ;
wire \bank_addr_this[1]~q ;
wire \row_mux_sel_last[1]~q ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \finished_tras_last~q ;
wire \p_main_fsm~171_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Selector42~7_combout ;
wire \Selector42~8_combout ;
wire \ba[1]~143_combout ;
wire \Selector10~2_combout ;
wire \writing_in_proc~2_combout ;
wire \writing_in_proc~q ;
wire \Selector5~4_combout ;
wire \Selector17~5_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \finished_tras~q ;
wire \p_main_fsm~161_combout ;
wire \p_main_fsm~164_combout ;
wire \p_main_fsm~165_combout ;
wire \Selector38~0_combout ;
wire \ba[1]~120_combout ;
wire \Selector42~5_combout ;
wire \Selector42~6_combout ;
wire \Selector2~14_combout ;
wire \Selector42~9_combout ;
wire \didnt_pch~q ;
wire \p_main_fsm~170_combout ;
wire \Selector5~6_combout ;
wire \Selector38~1_combout ;
wire \Selector38~2_combout ;
wire \didnt_act~q ;
wire \Selector10~1_combout ;
wire \Selector10~3_combout ;
wire \cs_n~64_combout ;
wire \Selector10~4_combout ;
wire \Selector10~5_combout ;
wire \state.s_holding~q ;
wire \Selector43~5_combout ;
wire \dqs_toggle_le_3~1_combout ;
wire \dqs_toggle_le_3~q ;
wire \Selector43~6_combout ;
wire \Selector43~7_combout ;
wire \Selector43~8_combout ;
wire \changing_cs_pause~q ;
wire \p_main_fsm~159_combout ;
wire \Selector12~6_combout ;
wire \Selector12~7_combout ;
wire \Selector12~8_combout ;
wire \state.s_writing~q ;
wire \wdata_burst_count[1]~50_combout ;
wire \Selector53~6_combout ;
wire \p_main_fsm~167_combout ;
wire \Selector53~8_combout ;
wire \wdata_burst_count[1]~68_combout ;
wire \Selector53~9_combout ;
wire \Selector53~10_combout ;
wire \Selector12~4_combout ;
wire \Selector46~14_combout ;
wire \Selector53~11_combout ;
wire \p_main_fsm~45_combout ;
wire \Selector0~19_combout ;
wire \Selector53~12_combout ;
wire \Selector53~13_combout ;
wire \Selector53~14_combout ;
wire \didnt_write~q ;
wire \Selector4~4_combout ;
wire \state.s_wait_for_init_done~1_combout ;
wire \state.s_wait_for_init_done~q ;
wire \Selector4~5_combout ;
wire \Selector4~6_combout ;
wire \Selector4~7_combout ;
wire \state.s_idle~q ;
wire \Selector20~19_combout ;
wire \Selector39~0_combout ;
wire \Selector39~1_combout ;
wire \Selector5~7_combout ;
wire \Selector39~2_combout ;
wire \doing_act~q ;
wire \trcd_pipe[0]~q ;
wire \finished_trcd~q ;
wire \ba[1]~123_combout ;
wire \Selector8~5_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \state.s_read~q ;
wire \Selector20~4_combout ;
wire \Selector46~8_combout ;
wire \new_req~45_combout ;
wire \new_req~46_combout ;
wire \new_req~47_combout ;
wire \Selector46~16_combout ;
wire \Selector46~9_combout ;
wire \Selector46~10_combout ;
wire \Selector46~11_combout ;
wire \process_13~0_combout ;
wire \Selector46~12_combout ;
wire \Selector46~13_combout ;
wire \new_req~q ;
wire \Selector11~1_combout ;
wire \new_req~49_combout ;
wire \Selector11~2_combout ;
wire \p_main_fsm~20_combout ;
wire \Selector11~4_combout ;
wire \Selector11~5_combout ;
wire \Selector11~6_combout ;
wire \state.s_reading~q ;
wire \ba[1]~119_combout ;
wire \Selector0~10_combout ;
wire \Selector0~11_combout ;
wire \Selector0~12_combout ;
wire \Selector0~17_combout ;
wire \Selector0~21_combout ;
wire \Selector0~22_combout ;
wire \Selector0~23_combout ;
wire \Selector0~4_combout ;
wire \Selector0~25_combout ;
wire \Selector0~26_combout ;
wire \accepted~q ;
wire \read_req_this~q ;
wire \p_main_fsm~157_combout ;
wire \state~332_combout ;
wire \am_writing~24_combout ;
wire \Selector50~1_combout ;
wire \Selector50~2_combout ;
wire \Selector50~3_combout ;
wire \Selector50~4_combout ;
wire \Selector50~6_combout ;
wire \Selector50~7_combout ;
wire \Selector50~8_combout ;
wire \am_writing~q ;
wire \Selector3~4_combout ;
wire \dqs_toggle_eq_0~1_combout ;
wire \dqs_toggle_eq_0~q ;
wire \p_main_fsm~162_combout ;
wire \Equal19~0_combout ;
wire \finished_tras_all~q ;
wire \p_main_fsm~163_combout ;
wire \Selector23~3_combout ;
wire \Selector21~0_combout ;
wire \refresh_in_progress~q ;
wire \p_main_fsm~57_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Selector2~7_combout ;
wire \Selector2~8_combout ;
wire \Selector2~13_combout ;
wire \Selector2~9_combout ;
wire \Selector2~10_combout ;
wire \Selector2~11_combout ;
wire \doing_pch~q ;
wire \trp_pipe[0]~q ;
wire \finished_trp~q ;
wire \Selector5~2_combout ;
wire \Selector3~2_combout ;
wire \doing_rfsh~q ;
wire \trfc_pipe[0]~q ;
wire \trfc_pipe[1]~q ;
wire \trfc_pipe[2]~q ;
wire \trfc_pipe[3]~q ;
wire \trfc_pipe[4]~q ;
wire \trfc_pipe[5]~q ;
wire \trfc_pipe[6]~q ;
wire \trfc_pipe[7]~q ;
wire \finished_trfc~q ;
wire \Selector3~3_combout ;
wire \state.s_refresh~q ;
wire \Selector2~12_combout ;
wire \state.s_precharge~q ;
wire \ba[1]~116_combout ;
wire \Selector15~0_combout ;
wire \rfsh_done~q ;
wire \rdata_valid_pipe~2_combout ;
wire \rdata_valid_pipe[2]~q ;
wire \a[5]~576_combout ;
wire \new_req~48_combout ;
wire \Selector17~2_combout ;
wire \cs_n~61_combout ;
wire \cs_n~62_combout ;
wire \Selector17~3_combout ;
wire \Selector17~6_combout ;
wire \Selector0~18_combout ;
wire \state~333_combout ;
wire \Selector17~8_combout ;
wire \p_main_fsm~169_combout ;
wire \Selector17~9_combout ;
wire \Selector17~10_combout ;
wire \Selector17~11_combout ;
wire \Selector17~12_combout ;
wire \Selector17~13_combout ;
wire \Selector17~15_combout ;
wire \Selector42~3_combout ;
wire \Selector17~16_combout ;
wire \Selector17~17_combout ;
wire \row_addr_this[0]~q ;
wire \a[0]~582_combout ;
wire \a[0]~583_combout ;
wire \a[5]~584_combout ;
wire \a[0]~585_combout ;
wire \a[0]~586_combout ;
wire \a[0]~587_combout ;
wire \Selector20~5_combout ;
wire \a[0]~588_combout ;
wire \a[0]~589_combout ;
wire \p_main_fsm~155_combout ;
wire \a[0]~590_combout ;
wire \Selector36~0_combout ;
wire \col_addr_next[0]~0_combout ;
wire \col_addr_this[0]~q ;
wire \row_addr_next[1]~1_combout ;
wire \row_addr_this[1]~q ;
wire \a[5]~594_combout ;
wire \a[5]~595_combout ;
wire \a[5]~597_combout ;
wire \a[5]~598_combout ;
wire \ba[1]~127_combout ;
wire \ba[1]~128_combout ;
wire \wdata_burst_count[1]~69_combout ;
wire \a[5]~599_combout ;
wire \a[5]~600_combout ;
wire \a[5]~605_combout ;
wire \a[5]~575_combout ;
wire \a[5]~606_combout ;
wire \a[5]~607_combout ;
wire \a[5]~596_combout ;
wire \a[5]~609_combout ;
wire \a[5]~610_combout ;
wire \a[5]~612_combout ;
wire \ba[1]~126_combout ;
wire \a[5]~592_combout ;
wire \a[5]~591_combout ;
wire \a[5]~613_combout ;
wire \a[5]~614_combout ;
wire \Selector35~0_combout ;
wire \col_addr_next[1]~1_combout ;
wire \col_addr_this[1]~q ;
wire \row_addr_this[2]~q ;
wire \Selector34~0_combout ;
wire \col_addr_next[2]~2_combout ;
wire \col_addr_this[2]~q ;
wire \row_addr_this[3]~q ;
wire \Selector33~0_combout ;
wire \col_addr_next[3]~3_combout ;
wire \col_addr_this[3]~q ;
wire \row_addr_next[4]~2_combout ;
wire \row_addr_this[4]~q ;
wire \Selector32~0_combout ;
wire \col_addr_next[4]~4_combout ;
wire \col_addr_this[4]~q ;
wire \row_addr_this[5]~q ;
wire \Selector31~0_combout ;
wire \col_addr_next[5]~5_combout ;
wire \col_addr_this[5]~q ;
wire \row_addr_next[6]~7_combout ;
wire \row_addr_this[6]~q ;
wire \Selector30~0_combout ;
wire \col_addr_next[6]~6_combout ;
wire \col_addr_this[6]~q ;
wire \row_addr_next[7]~8_combout ;
wire \row_addr_this[7]~q ;
wire \Selector29~0_combout ;
wire \col_addr_next[7]~7_combout ;
wire \col_addr_this[7]~q ;
wire \row_addr_this[8]~q ;
wire \Selector28~0_combout ;
wire \row_addr_next[9]~0_combout ;
wire \row_addr_this[9]~q ;
wire \Selector27~0_combout ;
wire \row_addr_next[10]~12_combout ;
wire \row_addr_this[10]~q ;
wire \Selector26~1_combout ;
wire \Selector26~2_combout ;
wire \Selector5~5_combout ;
wire \Selector26~0_combout ;
wire \Selector26~3_combout ;
wire \row_addr_this[11]~q ;
wire \Selector25~0_combout ;
wire \row_addr_this[12]~q ;
wire \Selector24~0_combout ;
wire \state~328_combout ;
wire \p_main_fsm~172_combout ;
wire \ba[1]~141_combout ;
wire \ba[1]~148_combout ;
wire \ba[1]~149_combout ;
wire \ba[1]~150_combout ;
wire \ba[1]~129_combout ;
wire \ba[1]~151_combout ;
wire \ba[1]~152_combout ;
wire \ba[1]~153_combout ;
wire \ba[1]~156_combout ;
wire \ba[1]~144_combout ;
wire \ba[1]~157_combout ;
wire \ba[1]~159_combout ;
wire \ba[1]~160_combout ;
wire \ba[1]~161_combout ;
wire \Selector41~0_combout ;
wire \Selector40~0_combout ;
wire \Selector18~0_combout ;
wire \Selector18~1_combout ;
wire \Selector18~3_combout ;
wire \Selector18~4_combout ;
wire \cs_n~63_combout ;
wire \Selector18~5_combout ;
wire \Selector18~6_combout ;
wire \Selector19~7_combout ;
wire \Selector12~2_combout ;
wire \Selector17~14_combout ;
wire \Selector19~10_combout ;
wire \p_main_fsm~168_combout ;
wire \Selector6~0_combout ;
wire \Selector19~8_combout ;
wire \Selector20~10_combout ;
wire \Selector20~11_combout ;
wire \Selector37~3_combout ;
wire \Selector20~12_combout ;
wire \Selector20~13_combout ;
wire \Selector20~14_combout ;
wire \Selector20~15_combout ;
wire \Selector20~16_combout ;
wire \p_main_fsm~173_combout ;
wire \Selector20~17_combout ;
wire \control_wlat_r[0]~0_combout ;
wire \control_wlat_r[1]~q ;
wire \control_wlat_r[4]~q ;
wire \control_wlat_r[3]~q ;
wire \control_wlat_r[2]~1_combout ;
wire \control_wlat_r[2]~q ;
wire \fifo_rdreq_cas4~q ;
wire \fifo_rdreq_cas5~q ;
wire \control_doing_wr~2_combout ;
wire \fifo_rdreq_cas6~q ;
wire \LessThan6~0_combout ;
wire \dqs_brst_odd_dtt~q ;


altera_ddr_auk_ddr_hp_avalon_if \g_local_avalon_if:av_if (
	.pipefull_3(\in_buf|my_fifo|pipefull[3]~q ),
	.clk(clk),
	.local_be({q_b_35,q_b_34,q_b_33,q_b_32}),
	.local_wdata({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.reset_phy_clk_1x_n(reset_n),
	.control_doing_wr(control_doing_wr1),
	.control_doing_wr1(control_doing_wr2),
	.local_write_req(local_write_req),
	.avalon_be({local_be_3,local_be_2,local_be_1,local_be_0}),
	.avalon_wdata({local_wdata_31,local_wdata_30,local_wdata_29,local_wdata_28,local_wdata_27,local_wdata_26,local_wdata_25,local_wdata_24,local_wdata_23,local_wdata_22,local_wdata_21,local_wdata_20,local_wdata_19,local_wdata_18,local_wdata_17,local_wdata_16,local_wdata_15,local_wdata_14,
local_wdata_13,local_wdata_12,local_wdata_11,local_wdata_10,local_wdata_9,local_wdata_8,local_wdata_7,local_wdata_6,local_wdata_5,local_wdata_4,local_wdata_3,local_wdata_2,local_wdata_1,local_wdata_0}));

altera_ddr_auk_ddr_hp_input_buf in_buf(
	.pipefull_3(\in_buf|my_fifo|pipefull[3]~q ),
	.clk(clk),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ready(ready1),
	.reset_n(reset_n),
	.write_req(\write_req_to_in_buf~0_combout ),
	.accepted(\accepted~q ),
	.pipefull_0(\in_buf|my_fifo|pipefull[0]~q ),
	.pipe_29_0(\in_buf|my_fifo|pipe[0][29]~q ),
	.pipe_28_0(\in_buf|my_fifo|pipe[0][28]~q ),
	.pipe_27_0(\in_buf|my_fifo|pipe[0][27]~q ),
	.pipe_9_0(\in_buf|my_fifo|pipe[0][9]~q ),
	.pipe_8_0(\in_buf|my_fifo|pipe[0][8]~q ),
	.pipe_19_0(\in_buf|my_fifo|pipe[0][19]~q ),
	.pipe_11_0(\in_buf|my_fifo|pipe[0][11]~q ),
	.pipe_14_0(\in_buf|my_fifo|pipe[0][14]~q ),
	.pipe_20_0(\in_buf|my_fifo|pipe[0][20]~q ),
	.pipe_18_0(\in_buf|my_fifo|pipe[0][18]~q ),
	.pipe_13_0(\in_buf|my_fifo|pipe[0][13]~q ),
	.pipe_15_0(\in_buf|my_fifo|pipe[0][15]~q ),
	.pipe_10_0(\in_buf|my_fifo|pipe[0][10]~q ),
	.pipe_16_0(\in_buf|my_fifo|pipe[0][16]~q ),
	.pipe_17_0(\in_buf|my_fifo|pipe[0][17]~q ),
	.pipe_21_0(\in_buf|my_fifo|pipe[0][21]~q ),
	.pipe_12_0(\in_buf|my_fifo|pipe[0][12]~q ),
	.pipe_22_0(\in_buf|my_fifo|pipe[0][22]~q ),
	.pipe_24_0(\in_buf|my_fifo|pipe[0][24]~q ),
	.pipe_25_0(\in_buf|my_fifo|pipe[0][25]~q ),
	.pipe_0_0(\in_buf|my_fifo|pipe[0][0]~q ),
	.pipe_1_0(\in_buf|my_fifo|pipe[0][1]~q ),
	.pipe_2_0(\in_buf|my_fifo|pipe[0][2]~q ),
	.pipe_3_0(\in_buf|my_fifo|pipe[0][3]~q ),
	.pipe_4_0(\in_buf|my_fifo|pipe[0][4]~q ),
	.pipe_5_0(\in_buf|my_fifo|pipe[0][5]~q ),
	.pipe_6_0(\in_buf|my_fifo|pipe[0][6]~q ),
	.pipe_7_0(\in_buf|my_fifo|pipe[0][7]~q ),
	.read_req(local_read_req),
	.row_addr({local_row_addr[12],local_row_addr[11],local_row_addr[10],local_row_addr[9],local_row_addr[8],local_row_addr[7],local_row_addr[6],local_row_addr[5],local_row_addr[4],local_row_addr[3],local_row_addr[2],local_row_addr[1],local_row_addr[0]}),
	.bank_addr({local_bank_addr[1],local_bank_addr[0]}),
	.size({local_size[1],local_size[0]}),
	.col_addr({local_col_addr[7],local_col_addr[6],local_col_addr[5],local_col_addr[4],local_col_addr[3],local_col_addr[2],local_col_addr[1],local_col_addr[0]}));

altera_ddr_auk_ddr_hp_bank_details bank_man(
	.clk(clk),
	.reset_n(reset_n),
	.Equal8(\bank_man|Equal8~0_combout ),
	.doing_act(\doing_act~q ),
	.in_this_bank({gnd,\bank_addr_this[1]~q ,\bank_addr_this[0]~q }),
	.doing_pch_all(\doing_pch_all~q ),
	.doing_pch(\doing_pch~q ),
	.row_mux_sel_next_1(\row_mux_sel_next[1]~0_combout ),
	.row_mux_sel_next_0(\row_mux_sel_next[0]~1_combout ),
	.Mux11(\bank_man|Mux11~1_combout ),
	.Mux3(\bank_man|Mux3~1_combout ),
	.Mux8(\bank_man|Mux8~1_combout ),
	.Mux2(\bank_man|Mux2~1_combout ),
	.Mux9(\bank_man|Mux9~1_combout ),
	.Mux4(\bank_man|Mux4~1_combout ),
	.Mux12(\bank_man|Mux12~1_combout ),
	.Mux7(\bank_man|Mux7~1_combout ),
	.Mux5(\bank_man|Mux5~1_combout ),
	.Mux6(\bank_man|Mux6~1_combout ),
	.Mux10(\bank_man|Mux10~1_combout ),
	.Mux1(\bank_man|Mux1~1_combout ),
	.Mux0(\bank_man|Mux0~1_combout ),
	.Mux13(\bank_man|Mux13~1_combout ),
	.row_addr_this_0(\row_addr_this[0]~q ),
	.row_addr_this_1(\row_addr_this[1]~q ),
	.row_addr_this_2(\row_addr_this[2]~q ),
	.row_addr_this_3(\row_addr_this[3]~q ),
	.row_addr_this_4(\row_addr_this[4]~q ),
	.row_addr_this_5(\row_addr_this[5]~q ),
	.row_addr_this_6(\row_addr_this[6]~q ),
	.row_addr_this_7(\row_addr_this[7]~q ),
	.row_addr_this_8(\row_addr_this[8]~q ),
	.row_addr_this_9(\row_addr_this[9]~q ),
	.row_addr_this_10(\row_addr_this[10]~q ),
	.row_addr_this_11(\row_addr_this[11]~q ),
	.row_addr_this_12(\row_addr_this[12]~q ));

altera_ddr_auk_ddr_hp_timers \g_timers:0:bank_timer (
	.clk(clk),
	.reset_n(reset_n),
	.am_writing(\am_writing~q ),
	.doing_act(\doing_act~q ),
	.twr_pipe_2(\g_timers:0:bank_timer|twr_pipe[2]~q ),
	.to_this_bank_0(\to_this_bank[0]~q ),
	.finished_twr1(\g_timers:0:bank_timer|finished_twr~combout ),
	.finished_tras1(\g_timers:0:bank_timer|finished_tras~q ));

altera_ddr_auk_ddr_hp_timers_1 \g_timers:1:bank_timer (
	.clk(clk),
	.reset_n(reset_n),
	.am_writing(\am_writing~q ),
	.doing_act(\doing_act~q ),
	.twr_pipe_2(\g_timers:1:bank_timer|twr_pipe[2]~q ),
	.to_this_bank_1(\to_this_bank[1]~q ),
	.finished_twr1(\g_timers:1:bank_timer|finished_twr~combout ),
	.finished_tras1(\g_timers:1:bank_timer|finished_tras~q ));

altera_ddr_auk_ddr_hp_timers_2 \g_timers:2:bank_timer (
	.clk(clk),
	.reset_n(reset_n),
	.am_writing(\am_writing~q ),
	.doing_act(\doing_act~q ),
	.twr_pipe_2(\g_timers:2:bank_timer|twr_pipe[2]~q ),
	.to_this_bank_2(\to_this_bank[2]~q ),
	.finished_twr1(\g_timers:2:bank_timer|finished_twr~combout ),
	.finished_tras1(\g_timers:2:bank_timer|finished_tras~q ));

altera_ddr_auk_ddr_hp_timers_3 \g_timers:3:bank_timer (
	.clk(clk),
	.reset_n(reset_n),
	.am_writing(\am_writing~q ),
	.doing_act(\doing_act~q ),
	.twr_pipe_2(\g_timers:3:bank_timer|twr_pipe[2]~q ),
	.to_this_bank_3(\to_this_bank[3]~q ),
	.finished_twr1(\g_timers:3:bank_timer|finished_twr~combout ),
	.finished_tras1(\g_timers:3:bank_timer|finished_tras~q ));

dffeas \rfsh_counter[10] (
	.clk(clk),
	.d(\rfsh_counter[10]~68_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[10]~q ),
	.prn(vcc));
defparam \rfsh_counter[10] .is_wysiwyg = "true";
defparam \rfsh_counter[10] .power_up = "low";

dffeas \rfsh_counter[3] (
	.clk(clk),
	.d(\rfsh_counter[3]~54_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[3]~q ),
	.prn(vcc));
defparam \rfsh_counter[3] .is_wysiwyg = "true";
defparam \rfsh_counter[3] .power_up = "low";

dffeas \rfsh_counter[5] (
	.clk(clk),
	.d(\rfsh_counter[5]~58_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[5]~q ),
	.prn(vcc));
defparam \rfsh_counter[5] .is_wysiwyg = "true";
defparam \rfsh_counter[5] .power_up = "low";

dffeas \rfsh_counter[15] (
	.clk(clk),
	.d(\rfsh_counter[15]~78_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[15]~q ),
	.prn(vcc));
defparam \rfsh_counter[15] .is_wysiwyg = "true";
defparam \rfsh_counter[15] .power_up = "low";

dffeas \rfsh_counter[11] (
	.clk(clk),
	.d(\rfsh_counter[11]~70_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[11]~q ),
	.prn(vcc));
defparam \rfsh_counter[11] .is_wysiwyg = "true";
defparam \rfsh_counter[11] .power_up = "low";

cycloneiii_lcell_comb \rfsh_counter[3]~54 (
	.dataa(\rfsh_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[2]~53 ),
	.combout(\rfsh_counter[3]~54_combout ),
	.cout(\rfsh_counter[3]~55 ));
defparam \rfsh_counter[3]~54 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[3]~54 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[5]~58 (
	.dataa(\rfsh_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[4]~57 ),
	.combout(\rfsh_counter[5]~58_combout ),
	.cout(\rfsh_counter[5]~59 ));
defparam \rfsh_counter[5]~58 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[5]~58 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[10]~68 (
	.dataa(\rfsh_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[9]~67 ),
	.combout(\rfsh_counter[10]~68_combout ),
	.cout(\rfsh_counter[10]~69 ));
defparam \rfsh_counter[10]~68 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[10]~68 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[11]~70 (
	.dataa(\rfsh_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[10]~69 ),
	.combout(\rfsh_counter[11]~70_combout ),
	.cout(\rfsh_counter[11]~71 ));
defparam \rfsh_counter[11]~70 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[11]~70 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[14]~76 (
	.dataa(\rfsh_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[13]~75 ),
	.combout(\rfsh_counter[14]~76_combout ),
	.cout(\rfsh_counter[14]~77 ));
defparam \rfsh_counter[14]~76 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[14]~76 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[15]~78 (
	.dataa(\rfsh_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\rfsh_counter[14]~77 ),
	.combout(\rfsh_counter[15]~78_combout ),
	.cout());
defparam \rfsh_counter[15]~78 .lut_mask = 16'h5A5A;
defparam \rfsh_counter[15]~78 .sum_lutc_input = "cin";

dffeas held_burstbegin(
	.clk(clk),
	.d(\held_burstbegin~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\held_burstbegin~q ),
	.prn(vcc));
defparam held_burstbegin.is_wysiwyg = "true";
defparam held_burstbegin.power_up = "low";

cycloneiii_lcell_comb \write_req_to_in_buf~0 (
	.dataa(local_write_req),
	.datab(\held_burstbegin~q ),
	.datac(local_burstbegin),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_req_to_in_buf~0_combout ),
	.cout());
defparam \write_req_to_in_buf~0 .lut_mask = 16'hFEFE;
defparam \write_req_to_in_buf~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector23~2 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~154_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
defparam \Selector23~2 .lut_mask = 16'hEEEE;
defparam \Selector23~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \held_burstbegin~2 (
	.dataa(\held_burstbegin~q ),
	.datab(local_burstbegin),
	.datac(local_write_req),
	.datad(ready1),
	.cin(gnd),
	.combout(\held_burstbegin~2_combout ),
	.cout());
defparam \held_burstbegin~2 .lut_mask = 16'hACFF;
defparam \held_burstbegin~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~5 (
	.dataa(\state.s_write~q ),
	.datab(gnd),
	.datac(\read_req_this~q ),
	.datad(\p_main_fsm~105_combout ),
	.cin(gnd),
	.combout(\Selector0~5_combout ),
	.cout());
defparam \Selector0~5 .lut_mask = 16'hAFFF;
defparam \Selector0~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~6 (
	.dataa(\Selector0~5_combout ),
	.datab(\write_req_next~0_combout ),
	.datac(\size_this[0]~q ),
	.datad(\size_this[1]~q ),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
defparam \Selector0~6 .lut_mask = 16'hFEFF;
defparam \Selector0~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~117 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~39_combout ),
	.datac(\read_req_this~q ),
	.datad(\p_main_fsm~45_combout ),
	.cin(gnd),
	.combout(\ba[1]~117_combout ),
	.cout());
defparam \ba[1]~117 .lut_mask = 16'hACFF;
defparam \ba[1]~117 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~7 (
	.dataa(\in_buf|my_fifo|pipe[0][28]~q ),
	.datab(\in_buf|my_fifo|pipefull[0]~q ),
	.datac(\accepted~q ),
	.datad(\size_this[1]~q ),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
defparam \Selector0~7 .lut_mask = 16'hEFFF;
defparam \Selector0~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~8 (
	.dataa(\p_main_fsm~19_combout ),
	.datab(\read_req_next~0_combout ),
	.datac(\Selector0~7_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
defparam \Selector0~8 .lut_mask = 16'hFAFC;
defparam \Selector0~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~9 (
	.dataa(\Selector0~27_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\ba[1]~117_combout ),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
defparam \Selector0~9 .lut_mask = 16'hFFFE;
defparam \Selector0~9 .sum_lutc_input = "datac";

dffeas write_req_last(
	.clk(clk),
	.d(\state.s_write~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_req_last~2_combout ),
	.q(\write_req_last~q ),
	.prn(vcc));
defparam write_req_last.is_wysiwyg = "true";
defparam write_req_last.power_up = "low";

cycloneiii_lcell_comb \Selector0~13 (
	.dataa(\finished_twtr~q ),
	.datab(\write_req_last~q ),
	.datac(\write_req_next~0_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
defparam \Selector0~13 .lut_mask = 16'hBFFF;
defparam \Selector0~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~3 (
	.dataa(\state.s_activate~q ),
	.datab(\doing_act~q ),
	.datac(gnd),
	.datad(\finished_trcd~q ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
defparam \Selector5~3 .lut_mask = 16'hEEFF;
defparam \Selector5~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~14 (
	.dataa(\Selector0~4_combout ),
	.datab(\dqs_toggle_le_1~q ),
	.datac(\Selector5~3_combout ),
	.datad(\writing_in_proc~q ),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
defparam \Selector0~14 .lut_mask = 16'hFEFF;
defparam \Selector0~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\am_reading~q ),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
defparam \Selector0~15 .lut_mask = 16'h0FFF;
defparam \Selector0~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~16 (
	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~14_combout ),
	.datac(\trcd_pipe[0]~q ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
defparam \Selector0~16 .lut_mask = 16'hFFFE;
defparam \Selector0~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~20 (
	.dataa(\state.s_write~q ),
	.datab(\Selector0~18_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\new_req~q ),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
defparam \Selector0~20 .lut_mask = 16'hFEFF;
defparam \Selector0~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~24 (
	.dataa(ctl_init_success),
	.datab(\in_buf|my_fifo|pipefull[0]~q ),
	.datac(gnd),
	.datad(\state.s_wait_for_init_done~q ),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
defparam \Selector0~24 .lut_mask = 16'hEEFF;
defparam \Selector0~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~6 (
	.dataa(\state~328_combout ),
	.datab(\a[5]~575_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\bank_man|Equal8~0_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
defparam \Selector2~6 .lut_mask = 16'hFEFF;
defparam \Selector2~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~160 (
	.dataa(\writing_in_proc~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(seq_ac_add_1t_ac_lat_internal),
	.cin(gnd),
	.combout(\p_main_fsm~160_combout ),
	.cout());
defparam \p_main_fsm~160 .lut_mask = 16'hAAFF;
defparam \p_main_fsm~160 .sum_lutc_input = "datac";

dffeas \to_this_bank[2] (
	.clk(clk),
	.d(\Decoder1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\to_this_bank[2]~q ),
	.prn(vcc));
defparam \to_this_bank[2] .is_wysiwyg = "true";
defparam \to_this_bank[2] .power_up = "low";

dffeas \to_this_bank[1] (
	.clk(clk),
	.d(\Decoder1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\to_this_bank[1]~q ),
	.prn(vcc));
defparam \to_this_bank[1] .is_wysiwyg = "true";
defparam \to_this_bank[1] .power_up = "low";

dffeas \to_this_bank[0] (
	.clk(clk),
	.d(\Decoder1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\to_this_bank[0]~q ),
	.prn(vcc));
defparam \to_this_bank[0] .is_wysiwyg = "true";
defparam \to_this_bank[0] .power_up = "low";

dffeas \to_this_bank[3] (
	.clk(clk),
	.d(\Decoder1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\to_this_bank[3]~q ),
	.prn(vcc));
defparam \to_this_bank[3] .is_wysiwyg = "true";
defparam \to_this_bank[3] .power_up = "low";

cycloneiii_lcell_comb \state~329 (
	.dataa(\didnt_read~q ),
	.datab(\didnt_write~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~329_combout ),
	.cout());
defparam \state~329 .lut_mask = 16'hEEEE;
defparam \state~329 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~330 (
	.dataa(\didnt_term~q ),
	.datab(\p_main_fsm~166_combout ),
	.datac(\state~329_combout ),
	.datad(\rdata_bcount_eq_1~q ),
	.cin(gnd),
	.combout(\state~330_combout ),
	.cout());
defparam \state~330 .lut_mask = 16'hFEFF;
defparam \state~330 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\state.s_reading~q ),
	.datab(gnd),
	.datac(\ba[1]~118_combout ),
	.datad(\state~330_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hAFFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~1 (
	.dataa(\state.s_write~q ),
	.datab(\ba[1]~120_combout ),
	.datac(\Selector42~11_combout ),
	.datad(\didnt_pch~q ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hEFFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~2 (
	.dataa(\size_last[0]~q ),
	.datab(\size_last[1]~q ),
	.datac(\p_main_fsm~167_combout ),
	.datad(\p_main_fsm~157_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
defparam \Selector4~2 .lut_mask = 16'h8BFF;
defparam \Selector4~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~3 (
	.dataa(\Selector4~0_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\state.s_read~q ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
defparam \Selector4~3 .lut_mask = 16'hFFFE;
defparam \Selector4~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~331 (
	.dataa(\p_main_fsm~154_combout ),
	.datab(\p_main_fsm~163_combout ),
	.datac(\bank_man|Equal8~0_combout ),
	.datad(\p_main_fsm~155_combout ),
	.cin(gnd),
	.combout(\state~331_combout ),
	.cout());
defparam \state~331 .lut_mask = 16'hACFF;
defparam \state~331 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~0 (
	.dataa(\state.s_writing~q ),
	.datab(\wdata_burst_count[1]~50_combout ),
	.datac(\state.s_idle~q ),
	.datad(\p_main_fsm~19_combout ),
	.cin(gnd),
	.combout(\Selector50~0_combout ),
	.cout());
defparam \Selector50~0 .lut_mask = 16'hFEFF;
defparam \Selector50~0 .sum_lutc_input = "datac";

dffeas doing_pch_all(
	.clk(clk),
	.d(\Selector23~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_pch_all~q ),
	.prn(vcc));
defparam doing_pch_all.is_wysiwyg = "true";
defparam doing_pch_all.power_up = "low";

cycloneiii_lcell_comb \Equal2~0 (
	.dataa(\bank_man|Mux11~1_combout ),
	.datab(\bank_man|Mux3~1_combout ),
	.datac(\row_addr_next[9]~0_combout ),
	.datad(\row_addr_next[1]~1_combout ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h6996;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~1 (
	.dataa(gnd),
	.datab(\bank_man|Mux2~1_combout ),
	.datac(\in_buf|my_fifo|pipefull[0]~q ),
	.datad(\in_buf|my_fifo|pipe[0][20]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hC33C;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~2 (
	.dataa(\Equal2~0_combout ),
	.datab(\bank_man|Mux8~1_combout ),
	.datac(\row_addr_next[4]~2_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hBEFF;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~5 (
	.dataa(\bank_man|Mux5~1_combout ),
	.datab(\bank_man|Mux6~1_combout ),
	.datac(\row_addr_next[6]~7_combout ),
	.datad(\row_addr_next[7]~8_combout ),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
defparam \Equal2~5 .lut_mask = 16'h6996;
defparam \Equal2~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~3 (
	.dataa(\state.s_writing~q ),
	.datab(\write_req_this~q ),
	.datac(\p_main_fsm~159_combout ),
	.datad(\didnt_write~q ),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
defparam \Selector20~3 .lut_mask = 16'hBFFF;
defparam \Selector20~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~4 (
	.dataa(\Selector5~3_combout ),
	.datab(\Selector20~3_combout ),
	.datac(\p_main_fsm~158_combout ),
	.datad(\ba[1]~121_combout ),
	.cin(gnd),
	.combout(\Selector46~4_combout ),
	.cout());
defparam \Selector46~4 .lut_mask = 16'hFFFE;
defparam \Selector46~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~5 (
	.dataa(\state.s_reading~q ),
	.datab(\didnt_term~q ),
	.datac(\read_req_this~q ),
	.datad(\didnt_read~q ),
	.cin(gnd),
	.combout(\Selector46~5_combout ),
	.cout());
defparam \Selector46~5 .lut_mask = 16'hEFFF;
defparam \Selector46~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~6 (
	.dataa(\Selector46~5_combout ),
	.datab(\state.s_activate~q ),
	.datac(\new_req~49_combout ),
	.datad(\Selector12~2_combout ),
	.cin(gnd),
	.combout(\Selector46~6_combout ),
	.cout());
defparam \Selector46~6 .lut_mask = 16'hFFFE;
defparam \Selector46~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~7 (
	.dataa(\new_req~47_combout ),
	.datab(\Selector46~15_combout ),
	.datac(\Selector46~4_combout ),
	.datad(\Selector46~6_combout ),
	.cin(gnd),
	.combout(\Selector46~7_combout ),
	.cout());
defparam \Selector46~7 .lut_mask = 16'hFFFE;
defparam \Selector46~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~3 (
	.dataa(\Selector50~5_combout ),
	.datab(\ba[1]~123_combout ),
	.datac(\Selector8~5_combout ),
	.datad(\p_main_fsm~45_combout ),
	.cin(gnd),
	.combout(\Selector8~3_combout ),
	.cout());
defparam \Selector8~3 .lut_mask = 16'hFEFF;
defparam \Selector8~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdata_bcount_le_1~3 (
	.dataa(gnd),
	.datab(\rdata_burst_count[1]~q ),
	.datac(\rdata_burst_count[0]~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\rdata_bcount_le_1~3_combout ),
	.cout());
defparam \rdata_bcount_le_1~3 .lut_mask = 16'h3FFF;
defparam \rdata_bcount_le_1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~52 (
	.dataa(\size_this[0]~q ),
	.datab(\wdata_burst_count[0]~q ),
	.datac(\size_this[1]~q ),
	.datad(\wdata_burst_count[1]~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~52_combout ),
	.cout());
defparam \wdata_burst_count[1]~52 .lut_mask = 16'h6996;
defparam \wdata_burst_count[1]~52 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~55 (
	.dataa(\p_main_fsm~154_combout ),
	.datab(gnd),
	.datac(\state.s_idle~q ),
	.datad(\state.s_write~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~55_combout ),
	.cout());
defparam \wdata_burst_count[1]~55 .lut_mask = 16'hAFFF;
defparam \wdata_burst_count[1]~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~2 (
	.dataa(\bank_is_open~q ),
	.datab(\new_req~q ),
	.datac(\read_req_this~q ),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\Selector42~2_combout ),
	.cout());
defparam \Selector42~2 .lut_mask = 16'hFFFE;
defparam \Selector42~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~57 (
	.dataa(\wdata_burst_count[1]~55_combout ),
	.datab(\wdata_burst_count[1]~56_combout ),
	.datac(\state.s_activate~q ),
	.datad(\state.s_writing~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~57_combout ),
	.cout());
defparam \wdata_burst_count[1]~57 .lut_mask = 16'hBFFF;
defparam \wdata_burst_count[1]~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~58 (
	.dataa(\p_main_fsm~61_combout ),
	.datab(\wdata_burst_count[1]~51_combout ),
	.datac(\this_row_is_open~q ),
	.datad(\state.s_writing~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~58_combout ),
	.cout());
defparam \wdata_burst_count[1]~58 .lut_mask = 16'h8BFF;
defparam \wdata_burst_count[1]~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~59 (
	.dataa(\state.s_activate~q ),
	.datab(\Selector4~4_combout ),
	.datac(\state.s_idle~q ),
	.datad(\p_main_fsm~45_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~59_combout ),
	.cout());
defparam \wdata_burst_count[1]~59 .lut_mask = 16'hA3FF;
defparam \wdata_burst_count[1]~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~61 (
	.dataa(\wdata_burst_count[1]~54_combout ),
	.datab(\wdata_burst_count[1]~57_combout ),
	.datac(\wdata_burst_count[1]~58_combout ),
	.datad(\wdata_burst_count[1]~60_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~61_combout ),
	.cout());
defparam \wdata_burst_count[1]~61 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[1]~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~62 (
	.dataa(\wdata_burst_count[1]~q ),
	.datab(\wdata_burst_count[0]~q ),
	.datac(\wdata_burst_count[1]~52_combout ),
	.datad(\wdata_burst_count[1]~61_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~62_combout ),
	.cout());
defparam \wdata_burst_count[1]~62 .lut_mask = 16'hF9F6;
defparam \wdata_burst_count[1]~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~64 (
	.dataa(\state.s_activate~q ),
	.datab(\wdata_burst_count[1]~63_combout ),
	.datac(\wdata_burst_count[1]~50_combout ),
	.datad(\state.s_writing~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~64_combout ),
	.cout());
defparam \wdata_burst_count[1]~64 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[1]~64 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdata_bcount_eq_1~2 (
	.dataa(\rdata_bcount_eq_1~q ),
	.datab(\size_last[1]~q ),
	.datac(gnd),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\rdata_bcount_eq_1~2_combout ),
	.cout());
defparam \rdata_bcount_eq_1~2 .lut_mask = 16'hEEFF;
defparam \rdata_bcount_eq_1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~0 (
	.dataa(\state.s_reading~q ),
	.datab(\state~330_combout ),
	.datac(\Selector0~28_combout ),
	.datad(\ba[1]~119_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'hFEFF;
defparam \Selector11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdata_bcount_eq_0~3 (
	.dataa(\rdata_burst_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rdata_burst_count[1]~q ),
	.cin(gnd),
	.combout(\rdata_bcount_eq_0~3_combout ),
	.cout());
defparam \rdata_bcount_eq_0~3 .lut_mask = 16'hAAFF;
defparam \rdata_bcount_eq_0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~1 (
	.dataa(\read_req_this~q ),
	.datab(\didnt_read~q ),
	.datac(\state.s_reading~q ),
	.datad(\didnt_term~q ),
	.cin(gnd),
	.combout(\Selector43~1_combout ),
	.cout());
defparam \Selector43~1 .lut_mask = 16'hFEFF;
defparam \Selector43~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~2 (
	.dataa(\p_main_fsm~158_combout ),
	.datab(\a[5]~574_combout ),
	.datac(\p_main_fsm~168_combout ),
	.datad(\Selector43~1_combout ),
	.cin(gnd),
	.combout(\Selector43~2_combout ),
	.cout());
defparam \Selector43~2 .lut_mask = 16'hFFFE;
defparam \Selector43~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~0 (
	.dataa(\read_req_this~q ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\p_main_fsm~39_combout ),
	.datad(\p_main_fsm~166_combout ),
	.cin(gnd),
	.combout(\Selector45~0_combout ),
	.cout());
defparam \Selector45~0 .lut_mask = 16'hEFFF;
defparam \Selector45~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~1 (
	.dataa(\state.s_idle~q ),
	.datab(\Selector45~0_combout ),
	.datac(\read_req_this~q ),
	.datad(\a[5]~576_combout ),
	.cin(gnd),
	.combout(\Selector45~1_combout ),
	.cout());
defparam \Selector45~1 .lut_mask = 16'hEFFF;
defparam \Selector45~1 .sum_lutc_input = "datac";

dffeas dqs_toggle_le_2(
	.clk(clk),
	.d(\dqs_toggle_le_2~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_toggle_le_2~q ),
	.prn(vcc));
defparam dqs_toggle_le_2.is_wysiwyg = "true";
defparam dqs_toggle_le_2.power_up = "low";

cycloneiii_lcell_comb \Selector43~4 (
	.dataa(\state.s_writing~q ),
	.datab(\write_req_this~q ),
	.datac(\didnt_write~q ),
	.datad(\dqs_toggle_le_2~q ),
	.cin(gnd),
	.combout(\Selector43~4_combout ),
	.cout());
defparam \Selector43~4 .lut_mask = 16'hBFFF;
defparam \Selector43~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~4 (
	.dataa(\size_last[1]~q ),
	.datab(\this_row_is_open~q ),
	.datac(\bank_is_open~q ),
	.datad(\new_req~q ),
	.cin(gnd),
	.combout(\Selector44~4_combout ),
	.cout());
defparam \Selector44~4 .lut_mask = 16'hBFFF;
defparam \Selector44~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~5 (
	.dataa(\Selector44~4_combout ),
	.datab(\state.s_read~q ),
	.datac(\state.s_reading~q ),
	.datad(\wdata_burst_count[1]~50_combout ),
	.cin(gnd),
	.combout(\Selector44~5_combout ),
	.cout());
defparam \Selector44~5 .lut_mask = 16'h8BFF;
defparam \Selector44~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~6 (
	.dataa(\didnt_term~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\p_main_fsm~166_combout ),
	.datad(\p_main_fsm~169_combout ),
	.cin(gnd),
	.combout(\Selector44~6_combout ),
	.cout());
defparam \Selector44~6 .lut_mask = 16'h8DFF;
defparam \Selector44~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~7 (
	.dataa(\didnt_read~q ),
	.datab(\Selector44~5_combout ),
	.datac(\state.s_reading~q ),
	.datad(\Selector44~6_combout ),
	.cin(gnd),
	.combout(\Selector44~7_combout ),
	.cout());
defparam \Selector44~7 .lut_mask = 16'hFFFE;
defparam \Selector44~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~8 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_read~q ),
	.datac(gnd),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\Selector44~8_combout ),
	.cout());
defparam \Selector44~8 .lut_mask = 16'hEEFF;
defparam \Selector44~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~10 (
	.dataa(\p_main_fsm~166_combout ),
	.datab(\Selector46~14_combout ),
	.datac(\rdata_bcount_eq_1~q ),
	.datad(\didnt_write~q ),
	.cin(gnd),
	.combout(\Selector44~10_combout ),
	.cout());
defparam \Selector44~10 .lut_mask = 16'hEFFF;
defparam \Selector44~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~3 (
	.dataa(\p_main_fsm~45_combout ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\Selector20~19_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
defparam \Selector12~3 .lut_mask = 16'hFEFF;
defparam \Selector12~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~5 (
	.dataa(\p_main_fsm~156_combout ),
	.datab(\Selector12~3_combout ),
	.datac(\Selector20~2_combout ),
	.datad(\Selector12~4_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
defparam \Selector12~5 .lut_mask = 16'hFFFE;
defparam \Selector12~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~7 (
	.dataa(\state.s_read~q ),
	.datab(\size_last[1]~q ),
	.datac(\state.s_writing~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector53~7_combout ),
	.cout());
defparam \Selector53~7 .lut_mask = 16'hFEFE;
defparam \Selector53~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \cs_n~60 (
	.dataa(\am_writing~q ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\cs_n~60_combout ),
	.cout());
defparam \cs_n~60 .lut_mask = 16'hAFFF;
defparam \cs_n~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~0 (
	.dataa(\cs_n~60_combout ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\cs_addr_to_term[0]~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'h8BFF;
defparam \Selector17~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~1 (
	.dataa(\Selector17~0_combout ),
	.datab(\a[5]~576_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector17~1_combout ),
	.cout());
defparam \Selector17~1 .lut_mask = 16'hEFFF;
defparam \Selector17~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~4 (
	.dataa(\p_main_fsm~165_combout ),
	.datab(gnd),
	.datac(\didnt_pch~q ),
	.datad(\didnt_act~q ),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
defparam \Selector17~4 .lut_mask = 16'hAFFF;
defparam \Selector17~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~7 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\size_last[1]~q ),
	.datad(\cs_addr_to_term[0]~q ),
	.cin(gnd),
	.combout(\Selector17~7_combout ),
	.cout());
defparam \Selector17~7 .lut_mask = 16'hACFF;
defparam \Selector17~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~577 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_write~q ),
	.datac(\state.s_read~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\a[0]~577_combout ),
	.cout());
defparam \a[0]~577 .lut_mask = 16'h8BFF;
defparam \a[0]~577 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~125 (
	.dataa(\state.s_precharge~q ),
	.datab(\finished_trp~q ),
	.datac(gnd),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\ba[1]~125_combout ),
	.cout());
defparam \ba[1]~125 .lut_mask = 16'hEEFF;
defparam \ba[1]~125 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~578 (
	.dataa(\state.s_precharge~q ),
	.datab(\a[0]~577_combout ),
	.datac(\ba[1]~125_combout ),
	.datad(\p_main_fsm~57_combout ),
	.cin(gnd),
	.combout(\a[0]~578_combout ),
	.cout());
defparam \a[0]~578 .lut_mask = 16'hFEFF;
defparam \a[0]~578 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~579 (
	.dataa(\state.s_read~q ),
	.datab(\bank_is_open~q ),
	.datac(\p_main_fsm~170_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[0]~579_combout ),
	.cout());
defparam \a[0]~579 .lut_mask = 16'hBFBF;
defparam \a[0]~579 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~580 (
	.dataa(\state.s_precharge~q ),
	.datab(\finished_trp~q ),
	.datac(\a[0]~579_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[0]~580_combout ),
	.cout());
defparam \a[0]~580 .lut_mask = 16'hD8D8;
defparam \a[0]~580 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~581 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_write~q ),
	.datac(\a[0]~580_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[0]~581_combout ),
	.cout());
defparam \a[0]~581 .lut_mask = 16'hFBFB;
defparam \a[0]~581 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~593 (
	.dataa(\Selector43~1_combout ),
	.datab(\a[5]~591_combout ),
	.datac(\p_main_fsm~158_combout ),
	.datad(\a[5]~592_combout ),
	.cin(gnd),
	.combout(\a[5]~593_combout ),
	.cout());
defparam \a[5]~593 .lut_mask = 16'hEFFF;
defparam \a[5]~593 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~601 (
	.dataa(\am_writing~q ),
	.datab(\state.s_idle~q ),
	.datac(\finished_trp~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\a[5]~601_combout ),
	.cout());
defparam \a[5]~601 .lut_mask = 16'h8BFF;
defparam \a[5]~601 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~602 (
	.dataa(\a[5]~601_combout ),
	.datab(\state.s_read~q ),
	.datac(\p_main_fsm~170_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\a[5]~602_combout ),
	.cout());
defparam \a[5]~602 .lut_mask = 16'hFEFF;
defparam \a[5]~602 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~603 (
	.dataa(\state.s_precharge~q ),
	.datab(\ba[1]~129_combout ),
	.datac(\p_main_fsm~57_combout ),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\a[5]~603_combout ),
	.cout());
defparam \a[5]~603 .lut_mask = 16'hEFFF;
defparam \a[5]~603 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~604 (
	.dataa(\a[5]~602_combout ),
	.datab(\a[5]~603_combout ),
	.datac(\a[5]~599_combout ),
	.datad(\a[5]~595_combout ),
	.cin(gnd),
	.combout(\a[5]~604_combout ),
	.cout());
defparam \a[5]~604 .lut_mask = 16'hFEFF;
defparam \a[5]~604 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~608 (
	.dataa(\state.s_reading~q ),
	.datab(\p_main_fsm~158_combout ),
	.datac(\a[5]~592_combout ),
	.datad(\ba[1]~118_combout ),
	.cin(gnd),
	.combout(\a[5]~608_combout ),
	.cout());
defparam \a[5]~608 .lut_mask = 16'hFEFF;
defparam \a[5]~608 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~611 (
	.dataa(\a[5]~584_combout ),
	.datab(\state~328_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\read_req_last~2_combout ),
	.cin(gnd),
	.combout(\a[5]~611_combout ),
	.cout());
defparam \a[5]~611 .lut_mask = 16'hFFEF;
defparam \a[5]~611 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~130 (
	.dataa(\state.s_precharge~q ),
	.datab(\state.s_idle~q ),
	.datac(\state.s_activate~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\ba[1]~130_combout ),
	.cout());
defparam \ba[1]~130 .lut_mask = 16'hFFFE;
defparam \ba[1]~130 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~131 (
	.dataa(\state.s_writing~q ),
	.datab(\p_main_fsm~159_combout ),
	.datac(\p_main_fsm~165_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ba[1]~131_combout ),
	.cout());
defparam \ba[1]~131 .lut_mask = 16'hB1B1;
defparam \ba[1]~131 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~132 (
	.dataa(\state.s_write~q ),
	.datab(\p_main_fsm~105_combout ),
	.datac(\ba[1]~130_combout ),
	.datad(\ba[1]~131_combout ),
	.cin(gnd),
	.combout(\ba[1]~132_combout ),
	.cout());
defparam \ba[1]~132 .lut_mask = 16'h27FF;
defparam \ba[1]~132 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~133 (
	.dataa(\state.s_read~q ),
	.datab(\state.s_precharge~q ),
	.datac(\state.s_idle~q ),
	.datad(\state.s_activate~q ),
	.cin(gnd),
	.combout(\ba[1]~133_combout ),
	.cout());
defparam \ba[1]~133 .lut_mask = 16'hBFFF;
defparam \ba[1]~133 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~134 (
	.dataa(\ba[1]~133_combout ),
	.datab(\cs_n~64_combout ),
	.datac(\finished_tras~q ),
	.datad(\finished_tras_last~q ),
	.cin(gnd),
	.combout(\ba[1]~134_combout ),
	.cout());
defparam \ba[1]~134 .lut_mask = 16'hFFFB;
defparam \ba[1]~134 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~135 (
	.dataa(\Mux2~1_combout ),
	.datab(\Mux3~1_combout ),
	.datac(\ba[1]~132_combout ),
	.datad(\ba[1]~134_combout ),
	.cin(gnd),
	.combout(\ba[1]~135_combout ),
	.cout());
defparam \ba[1]~135 .lut_mask = 16'hFFFE;
defparam \ba[1]~135 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~136 (
	.dataa(\state.s_read~q ),
	.datab(\state.s_precharge~q ),
	.datac(\state.s_activate~q ),
	.datad(\p_main_fsm~170_combout ),
	.cin(gnd),
	.combout(\ba[1]~136_combout ),
	.cout());
defparam \ba[1]~136 .lut_mask = 16'hBFFF;
defparam \ba[1]~136 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~137 (
	.dataa(\bank_is_open~q ),
	.datab(\state.s_idle~q ),
	.datac(\am_writing~q ),
	.datad(\ba[1]~136_combout ),
	.cin(gnd),
	.combout(\ba[1]~137_combout ),
	.cout());
defparam \ba[1]~137 .lut_mask = 16'hDF1F;
defparam \ba[1]~137 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~138 (
	.dataa(\p_main_fsm~63_combout ),
	.datab(\Selector50~5_combout ),
	.datac(gnd),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\ba[1]~138_combout ),
	.cout());
defparam \ba[1]~138 .lut_mask = 16'hAACC;
defparam \ba[1]~138 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~139 (
	.dataa(\ba[1]~125_combout ),
	.datab(\ba[1]~116_combout ),
	.datac(\state.s_activate~q ),
	.datad(\ba[1]~138_combout ),
	.cin(gnd),
	.combout(\ba[1]~139_combout ),
	.cout());
defparam \ba[1]~139 .lut_mask = 16'hFFFE;
defparam \ba[1]~139 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~140 (
	.dataa(\ba[1]~137_combout ),
	.datab(\ba[1]~139_combout ),
	.datac(\ba[1]~117_combout ),
	.datad(\p_main_fsm~156_combout ),
	.cin(gnd),
	.combout(\ba[1]~140_combout ),
	.cout());
defparam \ba[1]~140 .lut_mask = 16'hFFFE;
defparam \ba[1]~140 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~142 (
	.dataa(\state.s_precharge~q ),
	.datab(\state.s_holding~q ),
	.datac(gnd),
	.datad(\didnt_act~q ),
	.cin(gnd),
	.combout(\ba[1]~142_combout ),
	.cout());
defparam \ba[1]~142 .lut_mask = 16'hEEFF;
defparam \ba[1]~142 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_writing~q ),
	.datad(\didnt_pch~q ),
	.cin(gnd),
	.combout(\ba[1]~145_combout ),
	.cout());
defparam \ba[1]~145 .lut_mask = 16'h0FFF;
defparam \ba[1]~145 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~146 (
	.dataa(\wdata_burst_count[1]~51_combout ),
	.datab(\Selector4~4_combout ),
	.datac(\ba[1]~145_combout ),
	.datad(\state.s_precharge~q ),
	.cin(gnd),
	.combout(\ba[1]~146_combout ),
	.cout());
defparam \ba[1]~146 .lut_mask = 16'hFEFF;
defparam \ba[1]~146 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~147 (
	.dataa(\state.s_precharge~q ),
	.datab(\rfsh_pending~q ),
	.datac(\refresh_in_progress~q ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\ba[1]~147_combout ),
	.cout());
defparam \ba[1]~147 .lut_mask = 16'hFEFF;
defparam \ba[1]~147 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~154 (
	.dataa(\state.s_read~q ),
	.datab(\size_last[1]~q ),
	.datac(\write_req_this~q ),
	.datad(\ba[1]~121_combout ),
	.cin(gnd),
	.combout(\ba[1]~154_combout ),
	.cout());
defparam \ba[1]~154 .lut_mask = 16'hFFD8;
defparam \ba[1]~154 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~155 (
	.dataa(\ba[1]~124_combout ),
	.datab(\changing_cs_pause~q ),
	.datac(\p_main_fsm~155_combout ),
	.datad(\ba[1]~154_combout ),
	.cin(gnd),
	.combout(\ba[1]~155_combout ),
	.cout());
defparam \ba[1]~155 .lut_mask = 16'hFFEF;
defparam \ba[1]~155 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~158 (
	.dataa(\state.s_reading~q ),
	.datab(\p_main_fsm~158_combout ),
	.datac(\ba[1]~155_combout ),
	.datad(\ba[1]~118_combout ),
	.cin(gnd),
	.combout(\ba[1]~158_combout ),
	.cout());
defparam \ba[1]~158 .lut_mask = 16'hFEFF;
defparam \ba[1]~158 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~2 (
	.dataa(\am_writing~q ),
	.datab(\am_reading~q ),
	.datac(\finished_tras_all~q ),
	.datad(\this_row_is_open~q ),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
defparam \Selector18~2 .lut_mask = 16'hFFEF;
defparam \Selector18~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~6 (
	.dataa(\am_writing~q ),
	.datab(\am_reading~q ),
	.datac(\finished_tras_all~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
defparam \Selector20~6 .lut_mask = 16'hEFEF;
defparam \Selector20~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~7 (
	.dataa(\Selector20~19_combout ),
	.datab(\this_row_is_open~q ),
	.datac(\Selector20~2_combout ),
	.datad(\p_main_fsm~157_combout ),
	.cin(gnd),
	.combout(\Selector20~7_combout ),
	.cout());
defparam \Selector20~7 .lut_mask = 16'hFBFF;
defparam \Selector20~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~8 (
	.dataa(\Mux2~1_combout ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\Selector20~6_combout ),
	.datad(\Selector20~7_combout ),
	.cin(gnd),
	.combout(\Selector20~8_combout ),
	.cout());
defparam \Selector20~8 .lut_mask = 16'hFFF7;
defparam \Selector20~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~9 (
	.dataa(\this_row_is_open~q ),
	.datab(\Selector20~19_combout ),
	.datac(\read_req_this~q ),
	.datad(\p_main_fsm~45_combout ),
	.cin(gnd),
	.combout(\Selector20~9_combout ),
	.cout());
defparam \Selector20~9 .lut_mask = 16'hFFFE;
defparam \Selector20~9 .sum_lutc_input = "datac";

dffeas \bank_addr_this_valid[1] (
	.clk(clk),
	.d(\row_mux_sel_next[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_13~0_combout ),
	.q(\bank_addr_this_valid[1]~q ),
	.prn(vcc));
defparam \bank_addr_this_valid[1] .is_wysiwyg = "true";
defparam \bank_addr_this_valid[1] .power_up = "low";

dffeas \bank_addr_this_valid[0] (
	.clk(clk),
	.d(\row_mux_sel_next[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_13~0_combout ),
	.q(\bank_addr_this_valid[0]~q ),
	.prn(vcc));
defparam \bank_addr_this_valid[0] .is_wysiwyg = "true";
defparam \bank_addr_this_valid[0] .power_up = "low";

cycloneiii_lcell_comb \Decoder1~0 (
	.dataa(\bank_addr_this_valid[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\bank_addr_this_valid[0]~q ),
	.cin(gnd),
	.combout(\Decoder1~0_combout ),
	.cout());
defparam \Decoder1~0 .lut_mask = 16'hFF55;
defparam \Decoder1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Decoder1~1 (
	.dataa(\bank_addr_this_valid[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\bank_addr_this_valid[1]~q ),
	.cin(gnd),
	.combout(\Decoder1~1_combout ),
	.cout());
defparam \Decoder1~1 .lut_mask = 16'hFF55;
defparam \Decoder1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Decoder1~2 (
	.dataa(\bank_addr_this_valid[1]~q ),
	.datab(\bank_addr_this_valid[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder1~2_combout ),
	.cout());
defparam \Decoder1~2 .lut_mask = 16'hEEEE;
defparam \Decoder1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Decoder1~3 (
	.dataa(\bank_addr_this_valid[1]~q ),
	.datab(\bank_addr_this_valid[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder1~3_combout ),
	.cout());
defparam \Decoder1~3 .lut_mask = 16'h7777;
defparam \Decoder1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~18 (
	.dataa(\Selector20~19_combout ),
	.datab(\this_row_is_open~q ),
	.datac(\Mux2~1_combout ),
	.datad(\Selector20~6_combout ),
	.cin(gnd),
	.combout(\Selector20~18_combout ),
	.cout());
defparam \Selector20~18 .lut_mask = 16'hFFBF;
defparam \Selector20~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~4 (
	.dataa(\state~328_combout ),
	.datab(\Selector42~2_combout ),
	.datac(\Selector20~18_combout ),
	.datad(\Selector42~3_combout ),
	.cin(gnd),
	.combout(\Selector42~4_combout ),
	.cout());
defparam \Selector42~4 .lut_mask = 16'hFFFE;
defparam \Selector42~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~10 (
	.dataa(\state.s_write~q ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\state~328_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector42~10_combout ),
	.cout());
defparam \Selector42~10 .lut_mask = 16'hFEFF;
defparam \Selector42~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~0 (
	.dataa(\rfsh_counter[0]~q ),
	.datab(\rfsh_counter[1]~q ),
	.datac(\rfsh_counter[3]~q ),
	.datad(\rfsh_counter[4]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h7FFF;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~1 (
	.dataa(\rfsh_counter[11]~q ),
	.datab(\rfsh_counter[12]~q ),
	.datac(\rfsh_counter[13]~q ),
	.datad(\rfsh_counter[14]~q ),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~2 (
	.dataa(\rfsh_counter[10]~q ),
	.datab(\rfsh_counter[5]~q ),
	.datac(\rfsh_counter[6]~q ),
	.datad(\rfsh_counter[15]~q ),
	.cin(gnd),
	.combout(\LessThan0~2_combout ),
	.cout());
defparam \LessThan0~2 .lut_mask = 16'h7FFF;
defparam \LessThan0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~3 (
	.dataa(\rfsh_counter[2]~q ),
	.datab(\rfsh_counter[9]~q ),
	.datac(\rfsh_counter[7]~q ),
	.datad(\rfsh_counter[8]~q ),
	.cin(gnd),
	.combout(\LessThan0~3_combout ),
	.cout());
defparam \LessThan0~3 .lut_mask = 16'h7FFF;
defparam \LessThan0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan0~4 (
	.dataa(\LessThan0~0_combout ),
	.datab(\LessThan0~1_combout ),
	.datac(\LessThan0~2_combout ),
	.datad(\LessThan0~3_combout ),
	.cin(gnd),
	.combout(\LessThan0~4_combout ),
	.cout());
defparam \LessThan0~4 .lut_mask = 16'hFFFE;
defparam \LessThan0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[0]~70 (
	.dataa(\size_this[0]~q ),
	.datab(\wdata_burst_count[1]~q ),
	.datac(\wdata_burst_count[1]~61_combout ),
	.datad(\wdata_burst_count[0]~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[0]~70_combout ),
	.cout());
defparam \wdata_burst_count[0]~70 .lut_mask = 16'h6996;
defparam \wdata_burst_count[0]~70 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dqs_toggle_le_2~1 (
	.dataa(\state.s_write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\dqs_must_keep_toggling[2]~q ),
	.cin(gnd),
	.combout(\dqs_toggle_le_2~1_combout ),
	.cout());
defparam \dqs_toggle_le_2~1 .lut_mask = 16'hAAFF;
defparam \dqs_toggle_le_2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~27 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector0~27_combout ),
	.cout());
defparam \Selector0~27 .lut_mask = 16'hFFFE;
defparam \Selector0~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~11 (
	.dataa(\new_req~q ),
	.datab(\read_req_this~q ),
	.datac(\write_req_this~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector42~11_combout ),
	.cout());
defparam \Selector42~11 .lut_mask = 16'hFEFF;
defparam \Selector42~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~15 (
	.dataa(\size_last[1]~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\state.s_idle~q ),
	.datad(\new_req~48_combout ),
	.cin(gnd),
	.combout(\Selector46~15_combout ),
	.cout());
defparam \Selector46~15 .lut_mask = 16'hFFFD;
defparam \Selector46~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~9 (
	.dataa(\state.s_activate~q ),
	.datab(\finished_trcd~q ),
	.datac(\doing_act~q ),
	.datad(\Selector12~2_combout ),
	.cin(gnd),
	.combout(\Selector12~9_combout ),
	.cout());
defparam \Selector12~9 .lut_mask = 16'hFFEF;
defparam \Selector12~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~162 (
	.dataa(\state.s_holding~q ),
	.datab(\didnt_act~q ),
	.datac(\ba[1]~155_combout ),
	.datad(\a[5]~591_combout ),
	.cin(gnd),
	.combout(\ba[1]~162_combout ),
	.cout());
defparam \ba[1]~162 .lut_mask = 16'hFFFE;
defparam \ba[1]~162 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~9 (
	.dataa(\size_last[1]~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\new_req~48_combout ),
	.datad(\p_main_fsm~166_combout ),
	.cin(gnd),
	.combout(\Selector19~9_combout ),
	.cout());
defparam \Selector19~9 .lut_mask = 16'hFDFF;
defparam \Selector19~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb ready(
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(gnd),
	.datac(gnd),
	.datad(\in_buf|my_fifo|pipefull[3]~q ),
	.cin(gnd),
	.combout(ready1),
	.cout());
defparam ready.lut_mask = 16'hAAFF;
defparam ready.sum_lutc_input = "datac";

cycloneiii_lcell_comb local_refresh_ack(
	.dataa(ctl_init_success),
	.datab(\rfsh_done~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(local_refresh_ack1),
	.cout());
defparam local_refresh_ack.lut_mask = 16'hEEEE;
defparam local_refresh_ack.sum_lutc_input = "datac";

cycloneiii_lcell_comb \control_doing_rd[0] (
	.dataa(\state.s_read~q ),
	.datab(\rdata_valid_pipe[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(control_doing_rd_0),
	.cout());
defparam \control_doing_rd[0] .lut_mask = 16'hEEEE;
defparam \control_doing_rd[0] .sum_lutc_input = "datac";

dffeas \cs_n[0] (
	.clk(clk),
	.d(\Selector17~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cs_n_0),
	.prn(vcc));
defparam \cs_n[0] .is_wysiwyg = "true";
defparam \cs_n[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Selector36~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_0),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Selector35~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_1),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_2),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_3),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Selector32~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_4),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_5),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Selector30~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_6),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_7),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Selector28~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_8),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_9),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Selector26~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_10),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_11),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(a_12),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \ba[0] (
	.clk(clk),
	.d(\Selector41~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ba_0),
	.prn(vcc));
defparam \ba[0] .is_wysiwyg = "true";
defparam \ba[0] .power_up = "low";

dffeas \ba[1] (
	.clk(clk),
	.d(\Selector40~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ba_1),
	.prn(vcc));
defparam \ba[1] .is_wysiwyg = "true";
defparam \ba[1] .power_up = "low";

dffeas ras_n(
	.clk(clk),
	.d(\Selector18~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ras_n1),
	.prn(vcc));
defparam ras_n.is_wysiwyg = "true";
defparam ras_n.power_up = "low";

dffeas cas_n(
	.clk(clk),
	.d(\Selector19~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cas_n1),
	.prn(vcc));
defparam cas_n.is_wysiwyg = "true";
defparam cas_n.power_up = "low";

dffeas we_n(
	.clk(clk),
	.d(\Selector20~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(we_n1),
	.prn(vcc));
defparam we_n.is_wysiwyg = "true";
defparam we_n.power_up = "low";

dffeas \control_wlat_r[0] (
	.clk(clk),
	.d(\control_wlat_r[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(control_wlat_r_0),
	.prn(vcc));
defparam \control_wlat_r[0] .is_wysiwyg = "true";
defparam \control_wlat_r[0] .power_up = "low";

cycloneiii_lcell_comb \control_doing_wr~0 (
	.dataa(\control_wlat_r[1]~q ),
	.datab(\control_wlat_r[4]~q ),
	.datac(\control_wlat_r[3]~q ),
	.datad(\control_wlat_r[2]~q ),
	.cin(gnd),
	.combout(control_doing_wr),
	.cout());
defparam \control_doing_wr~0 .lut_mask = 16'hBFFF;
defparam \control_doing_wr~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal6~0 (
	.dataa(\control_wlat_r[1]~q ),
	.datab(\control_wlat_r[4]~q ),
	.datac(\control_wlat_r[3]~q ),
	.datad(\control_wlat_r[2]~q ),
	.cin(gnd),
	.combout(Equal6),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h7FFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \control_doing_wr~1 (
	.dataa(\fifo_rdreq_cas5~q ),
	.datab(control_wlat_r_0),
	.datac(control_doing_wr),
	.datad(Equal6),
	.cin(gnd),
	.combout(control_doing_wr1),
	.cout());
defparam \control_doing_wr~1 .lut_mask = 16'hBFFF;
defparam \control_doing_wr~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \control_doing_wr~3 (
	.dataa(\fifo_rdreq_cas4~q ),
	.datab(\control_doing_wr~2_combout ),
	.datac(\fifo_rdreq_cas6~q ),
	.datad(Equal6),
	.cin(gnd),
	.combout(control_doing_wr2),
	.cout());
defparam \control_doing_wr~3 .lut_mask = 16'hFAFC;
defparam \control_doing_wr~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \control_dqs_burst[0]~0 (
	.dataa(\dqs_must_keep_toggling[2]~q ),
	.datab(\dqs_must_keep_toggling[1]~q ),
	.datac(\dqs_must_keep_toggling[0]~q ),
	.datad(\dqs_brst_odd_dtt~q ),
	.cin(gnd),
	.combout(control_dqs_burst_0),
	.cout());
defparam \control_dqs_burst[0]~0 .lut_mask = 16'hFFFE;
defparam \control_dqs_burst[0]~0 .sum_lutc_input = "datac";

dffeas dqs_burst_cas4(
	.clk(clk),
	.d(dqs_burst_cas31),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_cas41),
	.prn(vcc));
defparam dqs_burst_cas4.is_wysiwyg = "true";
defparam dqs_burst_cas4.power_up = "low";

dffeas dqs_burst_cas3(
	.clk(clk),
	.d(control_dqs_burst_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_cas31),
	.prn(vcc));
defparam dqs_burst_cas3.is_wysiwyg = "true";
defparam dqs_burst_cas3.power_up = "low";

cycloneiii_lcell_comb \read_req_next~0 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_req_next~0_combout ),
	.cout());
defparam \read_req_next~0 .lut_mask = 16'hEEEE;
defparam \read_req_next~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rfsh_counter[0]~48 (
	.dataa(\LessThan0~4_combout ),
	.datab(\rfsh_counter[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\rfsh_counter[0]~48_combout ),
	.cout(\rfsh_counter[0]~49 ));
defparam \rfsh_counter[0]~48 .lut_mask = 16'h66EE;
defparam \rfsh_counter[0]~48 .sum_lutc_input = "datac";

dffeas \rfsh_counter[0] (
	.clk(clk),
	.d(\rfsh_counter[0]~48_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[0]~q ),
	.prn(vcc));
defparam \rfsh_counter[0] .is_wysiwyg = "true";
defparam \rfsh_counter[0] .power_up = "low";

cycloneiii_lcell_comb \rfsh_counter[1]~50 (
	.dataa(\rfsh_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[0]~49 ),
	.combout(\rfsh_counter[1]~50_combout ),
	.cout(\rfsh_counter[1]~51 ));
defparam \rfsh_counter[1]~50 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[1]~50 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[2]~52 (
	.dataa(\rfsh_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[1]~51 ),
	.combout(\rfsh_counter[2]~52_combout ),
	.cout(\rfsh_counter[2]~53 ));
defparam \rfsh_counter[2]~52 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[2]~52 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[4]~56 (
	.dataa(\rfsh_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[3]~55 ),
	.combout(\rfsh_counter[4]~56_combout ),
	.cout(\rfsh_counter[4]~57 ));
defparam \rfsh_counter[4]~56 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[4]~56 .sum_lutc_input = "cin";

dffeas \rfsh_counter[4] (
	.clk(clk),
	.d(\rfsh_counter[4]~56_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[4]~q ),
	.prn(vcc));
defparam \rfsh_counter[4] .is_wysiwyg = "true";
defparam \rfsh_counter[4] .power_up = "low";

dffeas \rfsh_counter[2] (
	.clk(clk),
	.d(\rfsh_counter[2]~52_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[2]~q ),
	.prn(vcc));
defparam \rfsh_counter[2] .is_wysiwyg = "true";
defparam \rfsh_counter[2] .power_up = "low";

dffeas \rfsh_counter[1] (
	.clk(clk),
	.d(\rfsh_counter[1]~50_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[1]~q ),
	.prn(vcc));
defparam \rfsh_counter[1] .is_wysiwyg = "true";
defparam \rfsh_counter[1] .power_up = "low";

cycloneiii_lcell_comb \LessThan1~0 (
	.dataa(\rfsh_counter[0]~q ),
	.datab(\rfsh_counter[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hEEEE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan1~1 (
	.dataa(\rfsh_counter[3]~q ),
	.datab(\rfsh_counter[4]~q ),
	.datac(\rfsh_counter[2]~q ),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hFFFE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rfsh_counter[6]~60 (
	.dataa(\rfsh_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[5]~59 ),
	.combout(\rfsh_counter[6]~60_combout ),
	.cout(\rfsh_counter[6]~61 ));
defparam \rfsh_counter[6]~60 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[6]~60 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[7]~62 (
	.dataa(\rfsh_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[6]~61 ),
	.combout(\rfsh_counter[7]~62_combout ),
	.cout(\rfsh_counter[7]~63 ));
defparam \rfsh_counter[7]~62 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[7]~62 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[8]~64 (
	.dataa(\rfsh_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[7]~63 ),
	.combout(\rfsh_counter[8]~64_combout ),
	.cout(\rfsh_counter[8]~65 ));
defparam \rfsh_counter[8]~64 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[8]~64 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \rfsh_counter[9]~66 (
	.dataa(\rfsh_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[8]~65 ),
	.combout(\rfsh_counter[9]~66_combout ),
	.cout(\rfsh_counter[9]~67 ));
defparam \rfsh_counter[9]~66 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[9]~66 .sum_lutc_input = "cin";

dffeas \rfsh_counter[9] (
	.clk(clk),
	.d(\rfsh_counter[9]~66_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[9]~q ),
	.prn(vcc));
defparam \rfsh_counter[9] .is_wysiwyg = "true";
defparam \rfsh_counter[9] .power_up = "low";

dffeas \rfsh_counter[6] (
	.clk(clk),
	.d(\rfsh_counter[6]~60_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[6]~q ),
	.prn(vcc));
defparam \rfsh_counter[6] .is_wysiwyg = "true";
defparam \rfsh_counter[6] .power_up = "low";

dffeas \rfsh_counter[7] (
	.clk(clk),
	.d(\rfsh_counter[7]~62_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[7]~q ),
	.prn(vcc));
defparam \rfsh_counter[7] .is_wysiwyg = "true";
defparam \rfsh_counter[7] .power_up = "low";

dffeas \rfsh_counter[8] (
	.clk(clk),
	.d(\rfsh_counter[8]~64_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[8]~q ),
	.prn(vcc));
defparam \rfsh_counter[8] .is_wysiwyg = "true";
defparam \rfsh_counter[8] .power_up = "low";

cycloneiii_lcell_comb \LessThan1~2 (
	.dataa(\rfsh_counter[5]~q ),
	.datab(\rfsh_counter[6]~q ),
	.datac(\rfsh_counter[7]~q ),
	.datad(\rfsh_counter[8]~q ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'hFFFE;
defparam \LessThan1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan1~3 (
	.dataa(\rfsh_counter[10]~q ),
	.datab(\LessThan1~1_combout ),
	.datac(\rfsh_counter[9]~q ),
	.datad(\LessThan1~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~3_combout ),
	.cout());
defparam \LessThan1~3 .lut_mask = 16'hFFFE;
defparam \LessThan1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rfsh_counter[12]~72 (
	.dataa(\rfsh_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[11]~71 ),
	.combout(\rfsh_counter[12]~72_combout ),
	.cout(\rfsh_counter[12]~73 ));
defparam \rfsh_counter[12]~72 .lut_mask = 16'h5AAF;
defparam \rfsh_counter[12]~72 .sum_lutc_input = "cin";

dffeas \rfsh_counter[12] (
	.clk(clk),
	.d(\rfsh_counter[12]~72_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[12]~q ),
	.prn(vcc));
defparam \rfsh_counter[12] .is_wysiwyg = "true";
defparam \rfsh_counter[12] .power_up = "low";

cycloneiii_lcell_comb \LessThan1~4 (
	.dataa(\rfsh_counter[11]~q ),
	.datab(\rfsh_counter[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~4_combout ),
	.cout());
defparam \LessThan1~4 .lut_mask = 16'hEEEE;
defparam \LessThan1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rfsh_counter[13]~74 (
	.dataa(\rfsh_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\rfsh_counter[12]~73 ),
	.combout(\rfsh_counter[13]~74_combout ),
	.cout(\rfsh_counter[13]~75 ));
defparam \rfsh_counter[13]~74 .lut_mask = 16'h5A5F;
defparam \rfsh_counter[13]~74 .sum_lutc_input = "cin";

dffeas \rfsh_counter[13] (
	.clk(clk),
	.d(\rfsh_counter[13]~74_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[13]~q ),
	.prn(vcc));
defparam \rfsh_counter[13] .is_wysiwyg = "true";
defparam \rfsh_counter[13] .power_up = "low";

dffeas \rfsh_counter[14] (
	.clk(clk),
	.d(\rfsh_counter[14]~76_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_counter[14]~q ),
	.prn(vcc));
defparam \rfsh_counter[14] .is_wysiwyg = "true";
defparam \rfsh_counter[14] .power_up = "low";

cycloneiii_lcell_comb \LessThan1~5 (
	.dataa(\rfsh_counter[15]~q ),
	.datab(\LessThan1~4_combout ),
	.datac(\rfsh_counter[13]~q ),
	.datad(\rfsh_counter[14]~q ),
	.cin(gnd),
	.combout(\LessThan1~5_combout ),
	.cout());
defparam \LessThan1~5 .lut_mask = 16'hFFFE;
defparam \LessThan1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rfsh_pending~2 (
	.dataa(\rfsh_pending~q ),
	.datab(ctl_init_success),
	.datac(\LessThan1~3_combout ),
	.datad(\LessThan1~5_combout ),
	.cin(gnd),
	.combout(\rfsh_pending~2_combout ),
	.cout());
defparam \rfsh_pending~2 .lut_mask = 16'hFFFE;
defparam \rfsh_pending~2 .sum_lutc_input = "datac";

dffeas rfsh_pending(
	.clk(clk),
	.d(\rfsh_pending~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\rfsh_done~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_pending~q ),
	.prn(vcc));
defparam rfsh_pending.is_wysiwyg = "true";
defparam rfsh_pending.power_up = "low";

cycloneiii_lcell_comb \size_next[1]~1 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\size_next[1]~1_combout ),
	.cout());
defparam \size_next[1]~1 .lut_mask = 16'hEEEE;
defparam \size_next[1]~1 .sum_lutc_input = "datac";

dffeas \size_this[1] (
	.clk(clk),
	.d(\size_next[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\size_this[1]~q ),
	.prn(vcc));
defparam \size_this[1] .is_wysiwyg = "true";
defparam \size_this[1] .power_up = "low";

dffeas accepted_r(
	.clk(clk),
	.d(\accepted~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\accepted_r~q ),
	.prn(vcc));
defparam accepted_r.is_wysiwyg = "true";
defparam accepted_r.power_up = "low";

dffeas \size_last[1] (
	.clk(clk),
	.d(\size_this[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\size_last[1]~q ),
	.prn(vcc));
defparam \size_last[1] .is_wysiwyg = "true";
defparam \size_last[1] .power_up = "low";

cycloneiii_lcell_comb \Selector37~2 (
	.dataa(\state.s_read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\size_last[1]~q ),
	.cin(gnd),
	.combout(\Selector37~2_combout ),
	.cout());
defparam \Selector37~2 .lut_mask = 16'hAAFF;
defparam \Selector37~2 .sum_lutc_input = "datac";

dffeas bank_is_open(
	.clk(clk),
	.d(\bank_man|Mux13~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bank_is_open~q ),
	.prn(vcc));
defparam bank_is_open.is_wysiwyg = "true";
defparam bank_is_open.power_up = "low";

cycloneiii_lcell_comb \size_next[0]~0 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\size_next[0]~0_combout ),
	.cout());
defparam \size_next[0]~0 .lut_mask = 16'hEEEE;
defparam \size_next[0]~0 .sum_lutc_input = "datac";

dffeas \size_this[0] (
	.clk(clk),
	.d(\size_next[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\size_this[0]~q ),
	.prn(vcc));
defparam \size_this[0] .is_wysiwyg = "true";
defparam \size_this[0] .power_up = "low";

dffeas \size_last[0] (
	.clk(clk),
	.d(\size_this[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted_r~q ),
	.q(\size_last[0]~q ),
	.prn(vcc));
defparam \size_last[0] .is_wysiwyg = "true";
defparam \size_last[0] .power_up = "low";

cycloneiii_lcell_comb \rdata_burst_count~6 (
	.dataa(\rdata_burst_count[1]~q ),
	.datab(\state.s_read~q ),
	.datac(\rdata_burst_count[0]~q ),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\rdata_burst_count~6_combout ),
	.cout());
defparam \rdata_burst_count~6 .lut_mask = 16'h8BFF;
defparam \rdata_burst_count~6 .sum_lutc_input = "datac";

dffeas \rdata_burst_count[0] (
	.clk(clk),
	.d(\rdata_burst_count~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_burst_count[0]~q ),
	.prn(vcc));
defparam \rdata_burst_count[0] .is_wysiwyg = "true";
defparam \rdata_burst_count[0] .power_up = "low";

cycloneiii_lcell_comb \rdata_burst_count~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\size_last[1]~q ),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\rdata_burst_count~4_combout ),
	.cout());
defparam \rdata_burst_count~4 .lut_mask = 16'h0FF0;
defparam \rdata_burst_count~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdata_burst_count~5 (
	.dataa(\rdata_burst_count[1]~q ),
	.datab(\rdata_burst_count[0]~q ),
	.datac(\state.s_read~q ),
	.datad(\rdata_burst_count~4_combout ),
	.cin(gnd),
	.combout(\rdata_burst_count~5_combout ),
	.cout());
defparam \rdata_burst_count~5 .lut_mask = 16'hACFF;
defparam \rdata_burst_count~5 .sum_lutc_input = "datac";

dffeas \rdata_burst_count[1] (
	.clk(clk),
	.d(\rdata_burst_count~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_burst_count[1]~q ),
	.prn(vcc));
defparam \rdata_burst_count[1] .is_wysiwyg = "true";
defparam \rdata_burst_count[1] .power_up = "low";

cycloneiii_lcell_comb \rdata_bcount_eq_1~3 (
	.dataa(\rdata_bcount_eq_1~2_combout ),
	.datab(\state.s_read~q ),
	.datac(\rdata_burst_count[1]~q ),
	.datad(\rdata_burst_count[0]~q ),
	.cin(gnd),
	.combout(\rdata_bcount_eq_1~3_combout ),
	.cout());
defparam \rdata_bcount_eq_1~3 .lut_mask = 16'hB8FF;
defparam \rdata_bcount_eq_1~3 .sum_lutc_input = "datac";

dffeas rdata_bcount_eq_1(
	.clk(clk),
	.d(\rdata_bcount_eq_1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_bcount_eq_1~q ),
	.prn(vcc));
defparam rdata_bcount_eq_1.is_wysiwyg = "true";
defparam rdata_bcount_eq_1.power_up = "low";

cycloneiii_lcell_comb \write_req_next~0 (
	.dataa(\in_buf|my_fifo|pipe[0][28]~q ),
	.datab(\in_buf|my_fifo|pipefull[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_req_next~0_combout ),
	.cout());
defparam \write_req_next~0 .lut_mask = 16'hEEEE;
defparam \write_req_next~0 .sum_lutc_input = "datac";

dffeas write_req_this(
	.clk(clk),
	.d(\write_req_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\write_req_this~q ),
	.prn(vcc));
defparam write_req_this.is_wysiwyg = "true";
defparam write_req_this.power_up = "low";

cycloneiii_lcell_comb \am_writing~25 (
	.dataa(\write_req_this~q ),
	.datab(\didnt_write~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\am_writing~25_combout ),
	.cout());
defparam \am_writing~25 .lut_mask = 16'hEEEE;
defparam \am_writing~25 .sum_lutc_input = "datac";

dffeas \rdata_valid_pipe[3] (
	.clk(clk),
	.d(control_doing_rd_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_valid_pipe[3]~q ),
	.prn(vcc));
defparam \rdata_valid_pipe[3] .is_wysiwyg = "true";
defparam \rdata_valid_pipe[3] .power_up = "low";

cycloneiii_lcell_comb \am_reading~0 (
	.dataa(\state.s_read~q ),
	.datab(\rdata_valid_pipe[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\am_reading~0_combout ),
	.cout());
defparam \am_reading~0 .lut_mask = 16'hEEEE;
defparam \am_reading~0 .sum_lutc_input = "datac";

dffeas am_reading(
	.clk(clk),
	.d(\am_reading~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\am_reading~q ),
	.prn(vcc));
defparam am_reading.is_wysiwyg = "true";
defparam am_reading.power_up = "low";

dffeas am_reading_r(
	.clk(clk),
	.d(\am_reading~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\am_reading_r~q ),
	.prn(vcc));
defparam am_reading_r.is_wysiwyg = "true";
defparam am_reading_r.power_up = "low";

cycloneiii_lcell_comb \Selector50~5 (
	.dataa(gnd),
	.datab(\am_writing~q ),
	.datac(\am_reading~q ),
	.datad(\am_reading_r~q ),
	.cin(gnd),
	.combout(\Selector50~5_combout ),
	.cout());
defparam \Selector50~5 .lut_mask = 16'h3FFF;
defparam \Selector50~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~105 (
	.dataa(\am_reading~q ),
	.datab(\size_last[1]~q ),
	.datac(gnd),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~105_combout ),
	.cout());
defparam \p_main_fsm~105 .lut_mask = 16'hEEFF;
defparam \p_main_fsm~105 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~8 (
	.dataa(\state.s_activate~q ),
	.datab(\doing_act~q ),
	.datac(\finished_trcd~q ),
	.datad(\Selector39~2_combout ),
	.cin(gnd),
	.combout(\Selector5~8_combout ),
	.cout());
defparam \Selector5~8 .lut_mask = 16'hFFEF;
defparam \Selector5~8 .sum_lutc_input = "datac";

dffeas \state.s_activate (
	.clk(clk),
	.d(\Selector5~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_activate~q ),
	.prn(vcc));
defparam \state.s_activate .is_wysiwyg = "true";
defparam \state.s_activate .power_up = "low";

cycloneiii_lcell_comb \wdata_burst_count[1]~53 (
	.dataa(\p_main_fsm~159_combout ),
	.datab(\state.s_writing~q ),
	.datac(\p_main_fsm~105_combout ),
	.datad(\state.s_activate~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~53_combout ),
	.cout());
defparam \wdata_burst_count[1]~53 .lut_mask = 16'h8BFF;
defparam \wdata_burst_count[1]~53 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~54 (
	.dataa(\state.s_activate~q ),
	.datab(\Selector50~5_combout ),
	.datac(\state.s_idle~q ),
	.datad(\wdata_burst_count[1]~53_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~54_combout ),
	.cout());
defparam \wdata_burst_count[1]~54 .lut_mask = 16'h7FFF;
defparam \wdata_burst_count[1]~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[8]~3 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[8]~3_combout ),
	.cout());
defparam \row_addr_next[8]~3 .lut_mask = 16'hEEEE;
defparam \row_addr_next[8]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[3]~4 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[3]~4_combout ),
	.cout());
defparam \row_addr_next[3]~4 .lut_mask = 16'hEEEE;
defparam \row_addr_next[3]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~3 (
	.dataa(\bank_man|Mux9~1_combout ),
	.datab(\bank_man|Mux4~1_combout ),
	.datac(\row_addr_next[8]~3_combout ),
	.datad(\row_addr_next[3]~4_combout ),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
defparam \Equal2~3 .lut_mask = 16'h6996;
defparam \Equal2~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[5]~5 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[5]~5_combout ),
	.cout());
defparam \row_addr_next[5]~5 .lut_mask = 16'hEEEE;
defparam \row_addr_next[5]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[0]~6 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[0]~6_combout ),
	.cout());
defparam \row_addr_next[0]~6 .lut_mask = 16'hEEEE;
defparam \row_addr_next[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~4 (
	.dataa(\bank_man|Mux12~1_combout ),
	.datab(\bank_man|Mux7~1_combout ),
	.datac(\row_addr_next[5]~5_combout ),
	.datad(\row_addr_next[0]~6_combout ),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
defparam \Equal2~4 .lut_mask = 16'h6996;
defparam \Equal2~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[11]~9 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[11]~9_combout ),
	.cout());
defparam \row_addr_next[11]~9 .lut_mask = 16'hEEEE;
defparam \row_addr_next[11]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[2]~10 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[2]~10_combout ),
	.cout());
defparam \row_addr_next[2]~10 .lut_mask = 16'hEEEE;
defparam \row_addr_next[2]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~6 (
	.dataa(\bank_man|Mux10~1_combout ),
	.datab(\bank_man|Mux1~1_combout ),
	.datac(\row_addr_next[11]~9_combout ),
	.datad(\row_addr_next[2]~10_combout ),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
defparam \Equal2~6 .lut_mask = 16'h6996;
defparam \Equal2~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[12]~11 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[12]~11_combout ),
	.cout());
defparam \row_addr_next[12]~11 .lut_mask = 16'hEEEE;
defparam \row_addr_next[12]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~7 (
	.dataa(\Equal2~5_combout ),
	.datab(\Equal2~6_combout ),
	.datac(\bank_man|Mux0~1_combout ),
	.datad(\row_addr_next[12]~11_combout ),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
defparam \Equal2~7 .lut_mask = 16'hEFFE;
defparam \Equal2~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal2~8 (
	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~3_combout ),
	.datac(\Equal2~4_combout ),
	.datad(\Equal2~7_combout ),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
defparam \Equal2~8 .lut_mask = 16'hFFFE;
defparam \Equal2~8 .sum_lutc_input = "datac";

dffeas this_row_is_open(
	.clk(clk),
	.d(\Equal2~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_buf|my_fifo|pipefull[0]~q ),
	.q(\this_row_is_open~q ),
	.prn(vcc));
defparam this_row_is_open.is_wysiwyg = "true";
defparam this_row_is_open.power_up = "low";

cycloneiii_lcell_comb \wdata_burst_count[1]~63 (
	.dataa(\wdata_burst_count[1]~51_combout ),
	.datab(\doing_act~q ),
	.datac(\finished_trcd~q ),
	.datad(\this_row_is_open~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~63_combout ),
	.cout());
defparam \wdata_burst_count[1]~63 .lut_mask = 16'h8DFF;
defparam \wdata_burst_count[1]~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~19 (
	.dataa(\size_last[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rdata_bcount_eq_1~q ),
	.cin(gnd),
	.combout(\p_main_fsm~19_combout ),
	.cout());
defparam \p_main_fsm~19 .lut_mask = 16'hAAFF;
defparam \p_main_fsm~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~2 (
	.dataa(\write_req_this~q ),
	.datab(\state.s_writing~q ),
	.datac(\p_main_fsm~159_combout ),
	.datad(\didnt_write~q ),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
defparam \Selector8~2 .lut_mask = 16'hFFFE;
defparam \Selector8~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~6 (
	.dataa(\p_main_fsm~105_combout ),
	.datab(\state.s_write~q ),
	.datac(\state~332_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(\Selector19~6_combout ),
	.cout());
defparam \Selector19~6 .lut_mask = 16'hBFFF;
defparam \Selector19~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~4 (
	.dataa(\Selector8~3_combout ),
	.datab(gnd),
	.datac(\read_req_this~q ),
	.datad(\Selector19~6_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
defparam \Selector8~4 .lut_mask = 16'hAFFF;
defparam \Selector8~4 .sum_lutc_input = "datac";

dffeas \state.s_write (
	.clk(clk),
	.d(\Selector8~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_write~q ),
	.prn(vcc));
defparam \state.s_write .is_wysiwyg = "true";
defparam \state.s_write .power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~154 (
	.dataa(\rfsh_pending~q ),
	.datab(\am_writing~q ),
	.datac(\am_reading~q ),
	.datad(\accepted_r~q ),
	.cin(gnd),
	.combout(\p_main_fsm~154_combout ),
	.cout());
defparam \p_main_fsm~154 .lut_mask = 16'hBFFF;
defparam \p_main_fsm~154 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~56 (
	.dataa(\Selector42~2_combout ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\state.s_write~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~56_combout ),
	.cout());
defparam \wdata_burst_count[1]~56 .lut_mask = 16'hACFF;
defparam \wdata_burst_count[1]~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~51 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_idle~q ),
	.datad(\state.s_write~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~51_combout ),
	.cout());
defparam \wdata_burst_count[1]~51 .lut_mask = 16'h0FFF;
defparam \wdata_burst_count[1]~51 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~65 (
	.dataa(\wdata_burst_count[1]~64_combout ),
	.datab(\wdata_burst_count[1]~63_combout ),
	.datac(\wdata_burst_count[1]~56_combout ),
	.datad(\wdata_burst_count[1]~51_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~65_combout ),
	.cout());
defparam \wdata_burst_count[1]~65 .lut_mask = 16'hEFFF;
defparam \wdata_burst_count[1]~65 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~122 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_idle~q ),
	.datad(\state.s_activate~q ),
	.cin(gnd),
	.combout(\ba[1]~122_combout ),
	.cout());
defparam \ba[1]~122 .lut_mask = 16'h0FFF;
defparam \ba[1]~122 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~60 (
	.dataa(\wdata_burst_count[1]~59_combout ),
	.datab(\state.s_writing~q ),
	.datac(\ba[1]~122_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~60_combout ),
	.cout());
defparam \wdata_burst_count[1]~60 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[1]~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~66 (
	.dataa(\Selector23~2_combout ),
	.datab(\wdata_burst_count[1]~54_combout ),
	.datac(\wdata_burst_count[1]~65_combout ),
	.datad(\wdata_burst_count[1]~60_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~66_combout ),
	.cout());
defparam \wdata_burst_count[1]~66 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[1]~66 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[0]~71 (
	.dataa(\wdata_burst_count[0]~70_combout ),
	.datab(\wdata_burst_count[1]~q ),
	.datac(\wdata_burst_count[0]~q ),
	.datad(\wdata_burst_count[1]~66_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[0]~71_combout ),
	.cout());
defparam \wdata_burst_count[0]~71 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[0]~71 .sum_lutc_input = "datac";

dffeas \wdata_burst_count[0] (
	.clk(clk),
	.d(\wdata_burst_count[0]~71_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_burst_count[0]~q ),
	.prn(vcc));
defparam \wdata_burst_count[0] .is_wysiwyg = "true";
defparam \wdata_burst_count[0] .power_up = "low";

cycloneiii_lcell_comb \wdata_burst_count[1]~67 (
	.dataa(\wdata_burst_count[1]~62_combout ),
	.datab(\wdata_burst_count[1]~q ),
	.datac(\wdata_burst_count[0]~q ),
	.datad(\wdata_burst_count[1]~66_combout ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~67_combout ),
	.cout());
defparam \wdata_burst_count[1]~67 .lut_mask = 16'hFEFF;
defparam \wdata_burst_count[1]~67 .sum_lutc_input = "datac";

dffeas \wdata_burst_count[1] (
	.clk(clk),
	.d(\wdata_burst_count[1]~67_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_burst_count[1]~q ),
	.prn(vcc));
defparam \wdata_burst_count[1] .is_wysiwyg = "true";
defparam \wdata_burst_count[1] .power_up = "low";

cycloneiii_lcell_comb \rdata_bcount_eq_0~4 (
	.dataa(\rdata_bcount_eq_0~3_combout ),
	.datab(\size_last[1]~q ),
	.datac(\rdata_bcount_eq_0~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\rdata_bcount_eq_0~4_combout ),
	.cout());
defparam \rdata_bcount_eq_0~4 .lut_mask = 16'hFFFD;
defparam \rdata_bcount_eq_0~4 .sum_lutc_input = "datac";

dffeas rdata_bcount_eq_0(
	.clk(clk),
	.d(\rdata_bcount_eq_0~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_bcount_eq_0~q ),
	.prn(vcc));
defparam rdata_bcount_eq_0.is_wysiwyg = "true";
defparam rdata_bcount_eq_0.power_up = "low";

dffeas \doing_wr_cl_pipe[0] (
	.clk(clk),
	.d(\am_writing~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_wr_cl_pipe[0]~q ),
	.prn(vcc));
defparam \doing_wr_cl_pipe[0] .is_wysiwyg = "true";
defparam \doing_wr_cl_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \finished_twtr~0 (
	.dataa(\am_writing~q ),
	.datab(\doing_wr_cl_pipe[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\finished_twtr~0_combout ),
	.cout());
defparam \finished_twtr~0 .lut_mask = 16'h7777;
defparam \finished_twtr~0 .sum_lutc_input = "datac";

dffeas finished_twtr(
	.clk(clk),
	.d(\finished_twtr~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_twtr~q ),
	.prn(vcc));
defparam finished_twtr.is_wysiwyg = "true";
defparam finished_twtr.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~158 (
	.dataa(\am_writing~q ),
	.datab(\rdata_bcount_eq_0~q ),
	.datac(\finished_twtr~q ),
	.datad(\changing_cs_pause~q ),
	.cin(gnd),
	.combout(\p_main_fsm~158_combout ),
	.cout());
defparam \p_main_fsm~158 .lut_mask = 16'hEFFF;
defparam \p_main_fsm~158 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dqs_must_keep_toggling[2]~8 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[1]~q ),
	.datac(\dqs_must_keep_toggling[0]~q ),
	.datad(\dqs_must_keep_toggling[2]~q ),
	.cin(gnd),
	.combout(\dqs_must_keep_toggling[2]~8_combout ),
	.cout());
defparam \dqs_must_keep_toggling[2]~8 .lut_mask = 16'hFFFD;
defparam \dqs_must_keep_toggling[2]~8 .sum_lutc_input = "datac";

dffeas \dqs_must_keep_toggling[2] (
	.clk(clk),
	.d(\dqs_must_keep_toggling[2]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_must_keep_toggling[2]~q ),
	.prn(vcc));
defparam \dqs_must_keep_toggling[2] .is_wysiwyg = "true";
defparam \dqs_must_keep_toggling[2] .power_up = "low";

cycloneiii_lcell_comb \dqs_must_keep_toggling[0]~7 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[0]~q ),
	.datac(\dqs_must_keep_toggling[2]~q ),
	.datad(\dqs_must_keep_toggling[1]~q ),
	.cin(gnd),
	.combout(\dqs_must_keep_toggling[0]~7_combout ),
	.cout());
defparam \dqs_must_keep_toggling[0]~7 .lut_mask = 16'hFFF7;
defparam \dqs_must_keep_toggling[0]~7 .sum_lutc_input = "datac";

dffeas \dqs_must_keep_toggling[0] (
	.clk(clk),
	.d(\dqs_must_keep_toggling[0]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_must_keep_toggling[0]~q ),
	.prn(vcc));
defparam \dqs_must_keep_toggling[0] .is_wysiwyg = "true";
defparam \dqs_must_keep_toggling[0] .power_up = "low";

cycloneiii_lcell_comb \dqs_must_keep_toggling[1]~6 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[1]~q ),
	.datac(\dqs_must_keep_toggling[0]~q ),
	.datad(\dqs_must_keep_toggling[2]~q ),
	.cin(gnd),
	.combout(\dqs_must_keep_toggling[1]~6_combout ),
	.cout());
defparam \dqs_must_keep_toggling[1]~6 .lut_mask = 16'hFFBE;
defparam \dqs_must_keep_toggling[1]~6 .sum_lutc_input = "datac";

dffeas \dqs_must_keep_toggling[1] (
	.clk(clk),
	.d(\dqs_must_keep_toggling[1]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_must_keep_toggling[1]~q ),
	.prn(vcc));
defparam \dqs_must_keep_toggling[1] .is_wysiwyg = "true";
defparam \dqs_must_keep_toggling[1] .power_up = "low";

cycloneiii_lcell_comb \dqs_toggle_le_1~1 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[1]~q ),
	.datac(\dqs_must_keep_toggling[0]~q ),
	.datad(\dqs_must_keep_toggling[2]~q ),
	.cin(gnd),
	.combout(\dqs_toggle_le_1~1_combout ),
	.cout());
defparam \dqs_toggle_le_1~1 .lut_mask = 16'hBFFF;
defparam \dqs_toggle_le_1~1 .sum_lutc_input = "datac";

dffeas dqs_toggle_le_1(
	.clk(clk),
	.d(\dqs_toggle_le_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_toggle_le_1~q ),
	.prn(vcc));
defparam dqs_toggle_le_1.is_wysiwyg = "true";
defparam dqs_toggle_le_1.power_up = "low";

cycloneiii_lcell_comb \Selector20~2 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_read~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector20~2_combout ),
	.cout());
defparam \Selector20~2 .lut_mask = 16'hEEEE;
defparam \Selector20~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rdata_bcount_le_1~4 (
	.dataa(\rdata_bcount_le_1~3_combout ),
	.datab(\size_last[0]~q ),
	.datac(\Selector20~2_combout ),
	.datad(\rdata_bcount_le_1~q ),
	.cin(gnd),
	.combout(\rdata_bcount_le_1~4_combout ),
	.cout());
defparam \rdata_bcount_le_1~4 .lut_mask = 16'hFFFD;
defparam \rdata_bcount_le_1~4 .sum_lutc_input = "datac";

dffeas rdata_bcount_le_1(
	.clk(clk),
	.d(\rdata_bcount_le_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_bcount_le_1~q ),
	.prn(vcc));
defparam rdata_bcount_le_1.is_wysiwyg = "true";
defparam rdata_bcount_le_1.power_up = "low";

cycloneiii_lcell_comb \a[5]~574 (
	.dataa(\finished_twtr~q ),
	.datab(\dqs_toggle_le_1~q ),
	.datac(gnd),
	.datad(\rdata_bcount_le_1~q ),
	.cin(gnd),
	.combout(\a[5]~574_combout ),
	.cout());
defparam \a[5]~574 .lut_mask = 16'hEEFF;
defparam \a[5]~574 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~166 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~166_combout ),
	.cout());
defparam \p_main_fsm~166 .lut_mask = 16'hFEFE;
defparam \p_main_fsm~166 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~3 (
	.dataa(\read_req_this~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
defparam \Selector11~3 .lut_mask = 16'hAAFF;
defparam \Selector11~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~39 (
	.dataa(\finished_twtr~q ),
	.datab(gnd),
	.datac(\am_writing~q ),
	.datad(\rdata_bcount_le_1~q ),
	.cin(gnd),
	.combout(\p_main_fsm~39_combout ),
	.cout());
defparam \p_main_fsm~39 .lut_mask = 16'hAFFF;
defparam \p_main_fsm~39 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~15 (
	.dataa(\state.s_idle~q ),
	.datab(\size_last[1]~q ),
	.datac(\rdata_bcount_eq_1~q ),
	.datad(\p_main_fsm~39_combout ),
	.cin(gnd),
	.combout(\Selector44~15_combout ),
	.cout());
defparam \Selector44~15 .lut_mask = 16'hEFFF;
defparam \Selector44~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~9 (
	.dataa(\Selector44~8_combout ),
	.datab(\Selector11~3_combout ),
	.datac(\state.s_write~q ),
	.datad(\Selector44~15_combout ),
	.cin(gnd),
	.combout(\Selector44~9_combout ),
	.cout());
defparam \Selector44~9 .lut_mask = 16'hFFFE;
defparam \Selector44~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~156 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~156_combout ),
	.cout());
defparam \p_main_fsm~156 .lut_mask = 16'hEEEE;
defparam \p_main_fsm~156 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~11 (
	.dataa(\accepted_r~q ),
	.datab(\p_main_fsm~156_combout ),
	.datac(\new_req~q ),
	.datad(\Selector37~2_combout ),
	.cin(gnd),
	.combout(\Selector44~11_combout ),
	.cout());
defparam \Selector44~11 .lut_mask = 16'hFFFE;
defparam \Selector44~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~63 (
	.dataa(\finished_twtr~q ),
	.datab(\dqs_toggle_le_1~q ),
	.datac(gnd),
	.datad(\rdata_bcount_eq_0~q ),
	.cin(gnd),
	.combout(\p_main_fsm~63_combout ),
	.cout());
defparam \p_main_fsm~63 .lut_mask = 16'hEEFF;
defparam \p_main_fsm~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~12 (
	.dataa(\Selector44~10_combout ),
	.datab(\Selector44~11_combout ),
	.datac(\ba[1]~123_combout ),
	.datad(\p_main_fsm~63_combout ),
	.cin(gnd),
	.combout(\Selector44~12_combout ),
	.cout());
defparam \Selector44~12 .lut_mask = 16'hFEFF;
defparam \Selector44~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~13 (
	.dataa(\read_req_this~q ),
	.datab(\p_main_fsm~166_combout ),
	.datac(\Selector44~9_combout ),
	.datad(\Selector44~12_combout ),
	.cin(gnd),
	.combout(\Selector44~13_combout ),
	.cout());
defparam \Selector44~13 .lut_mask = 16'hFFFE;
defparam \Selector44~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector37~6 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_read~q ),
	.datac(\state.s_reading~q ),
	.datad(\rdata_bcount_eq_1~q ),
	.cin(gnd),
	.combout(\Selector37~6_combout ),
	.cout());
defparam \Selector37~6 .lut_mask = 16'hFEFF;
defparam \Selector37~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~124 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_reading~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\ba[1]~124_combout ),
	.cout());
defparam \ba[1]~124 .lut_mask = 16'h0FFF;
defparam \ba[1]~124 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector37~4 (
	.dataa(\p_main_fsm~154_combout ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\ba[1]~124_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector37~4_combout ),
	.cout());
defparam \Selector37~4 .lut_mask = 16'hFAFC;
defparam \Selector37~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector37~5 (
	.dataa(\Selector37~3_combout ),
	.datab(\didnt_term~q ),
	.datac(\Selector37~6_combout ),
	.datad(\Selector37~4_combout ),
	.cin(gnd),
	.combout(\Selector37~5_combout ),
	.cout());
defparam \Selector37~5 .lut_mask = 16'hFFFE;
defparam \Selector37~5 .sum_lutc_input = "datac";

dffeas didnt_term(
	.clk(clk),
	.d(\Selector37~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\didnt_term~q ),
	.prn(vcc));
defparam didnt_term.is_wysiwyg = "true";
defparam didnt_term.power_up = "low";

cycloneiii_lcell_comb \Selector0~28 (
	.dataa(\read_req_this~q ),
	.datab(\didnt_read~q ),
	.datac(\didnt_term~q ),
	.datad(\p_main_fsm~158_combout ),
	.cin(gnd),
	.combout(\Selector0~28_combout ),
	.cout());
defparam \Selector0~28 .lut_mask = 16'hFFEF;
defparam \Selector0~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \read_req_last~3 (
	.dataa(\state.s_write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_req_last~3_combout ),
	.cout());
defparam \read_req_last~3 .lut_mask = 16'h5555;
defparam \read_req_last~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \read_req_last~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_write~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\read_req_last~2_combout ),
	.cout());
defparam \read_req_last~2 .lut_mask = 16'hFFF0;
defparam \read_req_last~2 .sum_lutc_input = "datac";

dffeas read_req_last(
	.clk(clk),
	.d(\read_req_last~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_req_last~2_combout ),
	.q(\read_req_last~q ),
	.prn(vcc));
defparam read_req_last.is_wysiwyg = "true";
defparam read_req_last.power_up = "low";

cycloneiii_lcell_comb \Selector45~2 (
	.dataa(\rdata_bcount_le_1~q ),
	.datab(\read_req_last~q ),
	.datac(\finished_twtr~q ),
	.datad(\dqs_toggle_le_1~q ),
	.cin(gnd),
	.combout(\Selector45~2_combout ),
	.cout());
defparam \Selector45~2 .lut_mask = 16'hEFFF;
defparam \Selector45~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~3 (
	.dataa(\state.s_reading~q ),
	.datab(\p_main_fsm~158_combout ),
	.datac(\Selector45~2_combout ),
	.datad(\ba[1]~118_combout ),
	.cin(gnd),
	.combout(\Selector45~3_combout ),
	.cout());
defparam \Selector45~3 .lut_mask = 16'hFEFF;
defparam \Selector45~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~61 (
	.dataa(\doing_act~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\finished_trcd~q ),
	.cin(gnd),
	.combout(\p_main_fsm~61_combout ),
	.cout());
defparam \p_main_fsm~61 .lut_mask = 16'hAAFF;
defparam \p_main_fsm~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~4 (
	.dataa(\state.s_activate~q ),
	.datab(\p_main_fsm~61_combout ),
	.datac(\read_req_this~q ),
	.datad(\p_main_fsm~63_combout ),
	.cin(gnd),
	.combout(\Selector45~4_combout ),
	.cout());
defparam \Selector45~4 .lut_mask = 16'hEFFF;
defparam \Selector45~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~5 (
	.dataa(\state.s_read~q ),
	.datab(\Selector45~4_combout ),
	.datac(\ba[1]~122_combout ),
	.datad(\state.s_reading~q ),
	.cin(gnd),
	.combout(\Selector45~5_combout ),
	.cout());
defparam \Selector45~5 .lut_mask = 16'hFEFF;
defparam \Selector45~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~6 (
	.dataa(\Selector45~1_combout ),
	.datab(\Selector45~3_combout ),
	.datac(\Selector45~5_combout ),
	.datad(\cs_addr_to_term[0]~q ),
	.cin(gnd),
	.combout(\Selector45~6_combout ),
	.cout());
defparam \Selector45~6 .lut_mask = 16'hFF7F;
defparam \Selector45~6 .sum_lutc_input = "datac";

dffeas \cs_addr_to_term[0] (
	.clk(clk),
	.d(\Selector45~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cs_addr_to_term[0]~q ),
	.prn(vcc));
defparam \cs_addr_to_term[0] .is_wysiwyg = "true";
defparam \cs_addr_to_term[0] .power_up = "low";

cycloneiii_lcell_comb \ba[1]~121 (
	.dataa(\state.s_reading~q ),
	.datab(\read_req_last~q ),
	.datac(\cs_addr_to_term[0]~q ),
	.datad(\a[5]~574_combout ),
	.cin(gnd),
	.combout(\ba[1]~121_combout ),
	.cout());
defparam \ba[1]~121 .lut_mask = 16'hEFFF;
defparam \ba[1]~121 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~14 (
	.dataa(\Selector44~7_combout ),
	.datab(\Selector44~13_combout ),
	.datac(\Selector0~28_combout ),
	.datad(\ba[1]~121_combout ),
	.cin(gnd),
	.combout(\Selector44~14_combout ),
	.cout());
defparam \Selector44~14 .lut_mask = 16'hFFFE;
defparam \Selector44~14 .sum_lutc_input = "datac";

dffeas didnt_read(
	.clk(clk),
	.d(\Selector44~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\didnt_read~q ),
	.prn(vcc));
defparam didnt_read.is_wysiwyg = "true";
defparam didnt_read.power_up = "low";

cycloneiii_lcell_comb \ba[1]~118 (
	.dataa(\read_req_this~q ),
	.datab(\didnt_read~q ),
	.datac(gnd),
	.datad(\didnt_term~q ),
	.cin(gnd),
	.combout(\ba[1]~118_combout ),
	.cout());
defparam \ba[1]~118 .lut_mask = 16'hEEFF;
defparam \ba[1]~118 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~3 (
	.dataa(\state.s_reading~q ),
	.datab(\p_main_fsm~158_combout ),
	.datac(\a[5]~574_combout ),
	.datad(\ba[1]~118_combout ),
	.cin(gnd),
	.combout(\Selector43~3_combout ),
	.cout());
defparam \Selector43~3 .lut_mask = 16'hEFFF;
defparam \Selector43~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_reading~q ),
	.datad(\state.s_writing~q ),
	.cin(gnd),
	.combout(\Selector43~0_combout ),
	.cout());
defparam \Selector43~0 .lut_mask = 16'h0FFF;
defparam \Selector43~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~0 (
	.dataa(\size_last[1]~q ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\state.s_read~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFEFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_mux_sel_next[0]~1 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_mux_sel_next[0]~1_combout ),
	.cout());
defparam \row_mux_sel_next[0]~1 .lut_mask = 16'hEEEE;
defparam \row_mux_sel_next[0]~1 .sum_lutc_input = "datac";

dffeas \bank_addr_this[0] (
	.clk(clk),
	.d(\row_mux_sel_next[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\bank_addr_this[0]~q ),
	.prn(vcc));
defparam \bank_addr_this[0] .is_wysiwyg = "true";
defparam \bank_addr_this[0] .power_up = "low";

cycloneiii_lcell_comb \row_mux_sel_next[1]~0 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_mux_sel_next[1]~0_combout ),
	.cout());
defparam \row_mux_sel_next[1]~0 .lut_mask = 16'hEEEE;
defparam \row_mux_sel_next[1]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_mux_sel_last[1]~2 (
	.dataa(\bank_addr_this[1]~q ),
	.datab(\row_mux_sel_next[1]~0_combout ),
	.datac(\bank_addr_this[0]~q ),
	.datad(\row_mux_sel_next[0]~1_combout ),
	.cin(gnd),
	.combout(\row_mux_sel_last[1]~2_combout ),
	.cout());
defparam \row_mux_sel_last[1]~2 .lut_mask = 16'h6996;
defparam \row_mux_sel_last[1]~2 .sum_lutc_input = "datac";

dffeas buf_not_empty_r(
	.clk(clk),
	.d(\in_buf|my_fifo|pipefull[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\buf_not_empty_r~q ),
	.prn(vcc));
defparam buf_not_empty_r.is_wysiwyg = "true";
defparam buf_not_empty_r.power_up = "low";

cycloneiii_lcell_comb \row_mux_sel_last[1]~3 (
	.dataa(\accepted_r~q ),
	.datab(\row_mux_sel_last[1]~2_combout ),
	.datac(\buf_not_empty_r~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_mux_sel_last[1]~3_combout ),
	.cout());
defparam \row_mux_sel_last[1]~3 .lut_mask = 16'hFEFE;
defparam \row_mux_sel_last[1]~3 .sum_lutc_input = "datac";

dffeas \row_mux_sel_last[0] (
	.clk(clk),
	.d(\bank_addr_this[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\row_mux_sel_last[1]~3_combout ),
	.q(\row_mux_sel_last[0]~q ),
	.prn(vcc));
defparam \row_mux_sel_last[0] .is_wysiwyg = "true";
defparam \row_mux_sel_last[0] .power_up = "low";

dffeas \bank_addr_this[1] (
	.clk(clk),
	.d(\row_mux_sel_next[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\bank_addr_this[1]~q ),
	.prn(vcc));
defparam \bank_addr_this[1] .is_wysiwyg = "true";
defparam \bank_addr_this[1] .power_up = "low";

dffeas \row_mux_sel_last[1] (
	.clk(clk),
	.d(\bank_addr_this[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\row_mux_sel_last[1]~3_combout ),
	.q(\row_mux_sel_last[1]~q ),
	.prn(vcc));
defparam \row_mux_sel_last[1] .is_wysiwyg = "true";
defparam \row_mux_sel_last[1] .power_up = "low";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(\row_mux_sel_last[0]~q ),
	.datab(\g_timers:2:bank_timer|finished_tras~q ),
	.datac(\row_mux_sel_last[1]~q ),
	.datad(\g_timers:0:bank_timer|finished_tras~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\g_timers:1:bank_timer|finished_tras~q ),
	.datab(\row_mux_sel_last[0]~q ),
	.datac(\Mux1~0_combout ),
	.datad(\g_timers:3:bank_timer|finished_tras~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

dffeas finished_tras_last(
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_tras_last~q ),
	.prn(vcc));
defparam finished_tras_last.is_wysiwyg = "true";
defparam finished_tras_last.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~171 (
	.dataa(\finished_tras~q ),
	.datab(\finished_tras_last~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~171_combout ),
	.cout());
defparam \p_main_fsm~171 .lut_mask = 16'hEEEE;
defparam \p_main_fsm~171 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(\row_mux_sel_last[1]~q ),
	.datab(\g_timers:1:bank_timer|finished_twr~combout ),
	.datac(\row_mux_sel_last[0]~q ),
	.datad(\g_timers:0:bank_timer|finished_twr~combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(\g_timers:2:bank_timer|finished_twr~combout ),
	.datab(\row_mux_sel_last[1]~q ),
	.datac(\Mux3~0_combout ),
	.datad(\g_timers:3:bank_timer|finished_twr~combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~7 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector42~7_combout ),
	.cout());
defparam \Selector42~7 .lut_mask = 16'hDDDD;
defparam \Selector42~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~8 (
	.dataa(\Mux2~1_combout ),
	.datab(\p_main_fsm~171_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\Selector42~7_combout ),
	.cin(gnd),
	.combout(\Selector42~8_combout ),
	.cout());
defparam \Selector42~8 .lut_mask = 16'hFF7F;
defparam \Selector42~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~143 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\ba[1]~143_combout ),
	.cout());
defparam \ba[1]~143 .lut_mask = 16'hFEFF;
defparam \ba[1]~143 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~2 (
	.dataa(\cs_n~62_combout ),
	.datab(\Selector10~0_combout ),
	.datac(\Selector42~8_combout ),
	.datad(\ba[1]~143_combout ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
defparam \Selector10~2 .lut_mask = 16'hFFFE;
defparam \Selector10~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \writing_in_proc~2 (
	.dataa(\writing_in_proc~q ),
	.datab(\state.s_write~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\writing_in_proc~2_combout ),
	.cout());
defparam \writing_in_proc~2 .lut_mask = 16'hEEEE;
defparam \writing_in_proc~2 .sum_lutc_input = "datac";

dffeas writing_in_proc(
	.clk(clk),
	.d(\writing_in_proc~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\am_writing~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\writing_in_proc~q ),
	.prn(vcc));
defparam writing_in_proc.is_wysiwyg = "true";
defparam writing_in_proc.power_up = "low";

cycloneiii_lcell_comb \Selector5~4 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\am_writing~q ),
	.datac(\writing_in_proc~q ),
	.datad(\changing_cs_pause~q ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
defparam \Selector5~4 .lut_mask = 16'hBFFF;
defparam \Selector5~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~5 (
	.dataa(\didnt_act~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector5~4_combout ),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
defparam \Selector17~5 .lut_mask = 16'hAAFF;
defparam \Selector17~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(\bank_addr_this[0]~q ),
	.datab(\g_timers:2:bank_timer|finished_tras~q ),
	.datac(\bank_addr_this[1]~q ),
	.datad(\g_timers:0:bank_timer|finished_tras~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(\g_timers:1:bank_timer|finished_tras~q ),
	.datab(\bank_addr_this[0]~q ),
	.datac(\Mux0~0_combout ),
	.datad(\g_timers:3:bank_timer|finished_tras~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

dffeas finished_tras(
	.clk(clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_tras~q ),
	.prn(vcc));
defparam finished_tras.is_wysiwyg = "true";
defparam finished_tras.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\am_writing~q ),
	.datad(\g_timers:2:bank_timer|twr_pipe[2]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~161_combout ),
	.cout());
defparam \p_main_fsm~161 .lut_mask = 16'h0FFF;
defparam \p_main_fsm~161 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~164 (
	.dataa(\finished_tras_last~q ),
	.datab(\g_timers:3:bank_timer|twr_pipe[2]~q ),
	.datac(\g_timers:1:bank_timer|twr_pipe[2]~q ),
	.datad(\g_timers:0:bank_timer|twr_pipe[2]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~164_combout ),
	.cout());
defparam \p_main_fsm~164 .lut_mask = 16'hFFFD;
defparam \p_main_fsm~164 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~165 (
	.dataa(\rdata_bcount_le_1~q ),
	.datab(\finished_tras~q ),
	.datac(\p_main_fsm~161_combout ),
	.datad(\p_main_fsm~164_combout ),
	.cin(gnd),
	.combout(\p_main_fsm~165_combout ),
	.cout());
defparam \p_main_fsm~165 .lut_mask = 16'hFFBF;
defparam \p_main_fsm~165 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector38~0 (
	.dataa(\state.s_read~q ),
	.datab(\state.s_holding~q ),
	.datac(\wdata_burst_count[1]~51_combout ),
	.datad(\Selector5~4_combout ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hBFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~120 (
	.dataa(\state.s_holding~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\didnt_act~q ),
	.cin(gnd),
	.combout(\ba[1]~120_combout ),
	.cout());
defparam \ba[1]~120 .lut_mask = 16'hAAFF;
defparam \ba[1]~120 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~5 (
	.dataa(gnd),
	.datab(\state.s_idle~q ),
	.datac(\state.s_write~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\Selector42~5_combout ),
	.cout());
defparam \Selector42~5 .lut_mask = 16'h3FFF;
defparam \Selector42~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~6 (
	.dataa(\didnt_pch~q ),
	.datab(\p_main_fsm~165_combout ),
	.datac(\ba[1]~120_combout ),
	.datad(\Selector42~5_combout ),
	.cin(gnd),
	.combout(\Selector42~6_combout ),
	.cout());
defparam \Selector42~6 .lut_mask = 16'hEFFF;
defparam \Selector42~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~14 (
	.dataa(\new_req~q ),
	.datab(\read_req_this~q ),
	.datac(\write_req_this~q ),
	.datad(\Selector20~2_combout ),
	.cin(gnd),
	.combout(\Selector2~14_combout ),
	.cout());
defparam \Selector2~14 .lut_mask = 16'hFFFE;
defparam \Selector2~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~9 (
	.dataa(\Selector42~4_combout ),
	.datab(\Selector42~6_combout ),
	.datac(\Selector2~14_combout ),
	.datad(\Selector42~8_combout ),
	.cin(gnd),
	.combout(\Selector42~9_combout ),
	.cout());
defparam \Selector42~9 .lut_mask = 16'hFFFE;
defparam \Selector42~9 .sum_lutc_input = "datac";

dffeas didnt_pch(
	.clk(clk),
	.d(\Selector42~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\didnt_pch~q ),
	.prn(vcc));
defparam didnt_pch.is_wysiwyg = "true";
defparam didnt_pch.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~170 (
	.dataa(\changing_cs_pause~q ),
	.datab(\didnt_pch~q ),
	.datac(\accepted_r~q ),
	.datad(seq_ac_add_1t_ac_lat_internal),
	.cin(gnd),
	.combout(\p_main_fsm~170_combout ),
	.cout());
defparam \p_main_fsm~170 .lut_mask = 16'hFEFF;
defparam \p_main_fsm~170 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~6 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(gnd),
	.datac(gnd),
	.datad(\am_writing~q ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
defparam \Selector5~6 .lut_mask = 16'hAAFF;
defparam \Selector5~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector38~1 (
	.dataa(\Selector2~14_combout ),
	.datab(\p_main_fsm~170_combout ),
	.datac(\ba[1]~143_combout ),
	.datad(\Selector5~6_combout ),
	.cin(gnd),
	.combout(\Selector38~1_combout ),
	.cout());
defparam \Selector38~1 .lut_mask = 16'hFEFF;
defparam \Selector38~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector38~2 (
	.dataa(\didnt_act~q ),
	.datab(\Selector38~0_combout ),
	.datac(\Selector38~1_combout ),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\Selector38~2_combout ),
	.cout());
defparam \Selector38~2 .lut_mask = 16'hFEFF;
defparam \Selector38~2 .sum_lutc_input = "datac";

dffeas didnt_act(
	.clk(clk),
	.d(\Selector38~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\didnt_act~q ),
	.prn(vcc));
defparam didnt_act.is_wysiwyg = "true";
defparam didnt_act.power_up = "low";

cycloneiii_lcell_comb \Selector10~1 (
	.dataa(\didnt_pch~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\didnt_act~q ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hAAFF;
defparam \Selector10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~3 (
	.dataa(\state.s_holding~q ),
	.datab(\Selector17~5_combout ),
	.datac(\p_main_fsm~165_combout ),
	.datad(\Selector10~1_combout ),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
defparam \Selector10~3 .lut_mask = 16'hFFFE;
defparam \Selector10~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \cs_n~64 (
	.dataa(\p_main_fsm~170_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\cs_n~64_combout ),
	.cout());
defparam \cs_n~64 .lut_mask = 16'hAAFF;
defparam \cs_n~64 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~4 (
	.dataa(\cs_n~60_combout ),
	.datab(\cs_n~64_combout ),
	.datac(\Selector10~0_combout ),
	.datad(\ba[1]~143_combout ),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
defparam \Selector10~4 .lut_mask = 16'hFFFE;
defparam \Selector10~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~5 (
	.dataa(\Selector42~10_combout ),
	.datab(\Selector10~2_combout ),
	.datac(\Selector10~3_combout ),
	.datad(\Selector10~4_combout ),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
defparam \Selector10~5 .lut_mask = 16'hFFFE;
defparam \Selector10~5 .sum_lutc_input = "datac";

dffeas \state.s_holding (
	.clk(clk),
	.d(\Selector10~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_holding~q ),
	.prn(vcc));
defparam \state.s_holding .is_wysiwyg = "true";
defparam \state.s_holding .power_up = "low";

cycloneiii_lcell_comb \Selector43~5 (
	.dataa(\Selector43~4_combout ),
	.datab(\Selector43~0_combout ),
	.datac(\state.s_idle~q ),
	.datad(\state.s_holding~q ),
	.cin(gnd),
	.combout(\Selector43~5_combout ),
	.cout());
defparam \Selector43~5 .lut_mask = 16'hEFFF;
defparam \Selector43~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dqs_toggle_le_3~1 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[2]~q ),
	.datac(\dqs_must_keep_toggling[1]~q ),
	.datad(\dqs_must_keep_toggling[0]~q ),
	.cin(gnd),
	.combout(\dqs_toggle_le_3~1_combout ),
	.cout());
defparam \dqs_toggle_le_3~1 .lut_mask = 16'hEFFF;
defparam \dqs_toggle_le_3~1 .sum_lutc_input = "datac";

dffeas dqs_toggle_le_3(
	.clk(clk),
	.d(\dqs_toggle_le_3~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_toggle_le_3~q ),
	.prn(vcc));
defparam dqs_toggle_le_3.is_wysiwyg = "true";
defparam dqs_toggle_le_3.power_up = "low";

cycloneiii_lcell_comb \Selector43~6 (
	.dataa(\state.s_holding~q ),
	.datab(\didnt_act~q ),
	.datac(\dqs_toggle_le_3~q ),
	.datad(\read_req_last~2_combout ),
	.cin(gnd),
	.combout(\Selector43~6_combout ),
	.cout());
defparam \Selector43~6 .lut_mask = 16'hFFBF;
defparam \Selector43~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~7 (
	.dataa(\Selector45~1_combout ),
	.datab(\Selector43~3_combout ),
	.datac(\Selector43~5_combout ),
	.datad(\Selector43~6_combout ),
	.cin(gnd),
	.combout(\Selector43~7_combout ),
	.cout());
defparam \Selector43~7 .lut_mask = 16'hFFFE;
defparam \Selector43~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~8 (
	.dataa(\Selector43~2_combout ),
	.datab(\changing_cs_pause~q ),
	.datac(\Selector43~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector43~8_combout ),
	.cout());
defparam \Selector43~8 .lut_mask = 16'hFEFE;
defparam \Selector43~8 .sum_lutc_input = "datac";

dffeas changing_cs_pause(
	.clk(clk),
	.d(\Selector43~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\changing_cs_pause~q ),
	.prn(vcc));
defparam changing_cs_pause.is_wysiwyg = "true";
defparam changing_cs_pause.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~159 (
	.dataa(\am_reading~q ),
	.datab(\am_reading_r~q ),
	.datac(\wdata_burst_count[1]~q ),
	.datad(\changing_cs_pause~q ),
	.cin(gnd),
	.combout(\p_main_fsm~159_combout ),
	.cout());
defparam \p_main_fsm~159 .lut_mask = 16'h7FFF;
defparam \p_main_fsm~159 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~6 (
	.dataa(\Selector12~9_combout ),
	.datab(\state.s_writing~q ),
	.datac(\am_writing~25_combout ),
	.datad(\p_main_fsm~159_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
defparam \Selector12~6 .lut_mask = 16'hFEFF;
defparam \Selector12~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~7 (
	.dataa(\state.s_write~q ),
	.datab(\am_reading~q ),
	.datac(\size_last[1]~q ),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\Selector12~7_combout ),
	.cout());
defparam \Selector12~7 .lut_mask = 16'hFEFF;
defparam \Selector12~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~8 (
	.dataa(\Selector12~5_combout ),
	.datab(\Selector12~6_combout ),
	.datac(\state~332_combout ),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector12~8_combout ),
	.cout());
defparam \Selector12~8 .lut_mask = 16'hFFFE;
defparam \Selector12~8 .sum_lutc_input = "datac";

dffeas \state.s_writing (
	.clk(clk),
	.d(\Selector12~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_writing~q ),
	.prn(vcc));
defparam \state.s_writing .is_wysiwyg = "true";
defparam \state.s_writing .power_up = "low";

cycloneiii_lcell_comb \wdata_burst_count[1]~50 (
	.dataa(gnd),
	.datab(\state.s_idle~q ),
	.datac(\state.s_write~q ),
	.datad(\state.s_activate~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~50_combout ),
	.cout());
defparam \wdata_burst_count[1]~50 .lut_mask = 16'h3FFF;
defparam \wdata_burst_count[1]~50 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~6 (
	.dataa(\write_req_this~q ),
	.datab(\state.s_writing~q ),
	.datac(\p_main_fsm~159_combout ),
	.datad(\wdata_burst_count[1]~50_combout ),
	.cin(gnd),
	.combout(\Selector53~6_combout ),
	.cout());
defparam \Selector53~6 .lut_mask = 16'hBFFF;
defparam \Selector53~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~167 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\new_req~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~167_combout ),
	.cout());
defparam \p_main_fsm~167 .lut_mask = 16'hFEFE;
defparam \p_main_fsm~167 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~8 (
	.dataa(\Selector53~7_combout ),
	.datab(\ba[1]~124_combout ),
	.datac(\p_main_fsm~167_combout ),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\Selector53~8_combout ),
	.cout());
defparam \Selector53~8 .lut_mask = 16'hEFFF;
defparam \Selector53~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~68 (
	.dataa(\read_req_this~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.s_writing~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~68_combout ),
	.cout());
defparam \wdata_burst_count[1]~68 .lut_mask = 16'hAAFF;
defparam \wdata_burst_count[1]~68 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~9 (
	.dataa(\state.s_reading~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\didnt_term~q ),
	.datad(\wdata_burst_count[1]~68_combout ),
	.cin(gnd),
	.combout(\Selector53~9_combout ),
	.cout());
defparam \Selector53~9 .lut_mask = 16'hEFFF;
defparam \Selector53~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~10 (
	.dataa(\didnt_write~q ),
	.datab(\Selector53~6_combout ),
	.datac(\Selector53~8_combout ),
	.datad(\Selector53~9_combout ),
	.cin(gnd),
	.combout(\Selector53~10_combout ),
	.cout());
defparam \Selector53~10 .lut_mask = 16'hFFFE;
defparam \Selector53~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~4 (
	.dataa(\new_req~q ),
	.datab(\write_req_this~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
defparam \Selector12~4 .lut_mask = 16'hEEEE;
defparam \Selector12~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~14 (
	.dataa(\didnt_term~q ),
	.datab(\state.s_reading~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector46~14_combout ),
	.cout());
defparam \Selector46~14 .lut_mask = 16'hEEEE;
defparam \Selector46~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~11 (
	.dataa(\state.s_read~q ),
	.datab(\Selector46~14_combout ),
	.datac(\rdata_bcount_eq_1~q ),
	.datad(\didnt_read~q ),
	.cin(gnd),
	.combout(\Selector53~11_combout ),
	.cout());
defparam \Selector53~11 .lut_mask = 16'hEFFF;
defparam \Selector53~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~45 (
	.dataa(\am_reading~q ),
	.datab(\am_reading_r~q ),
	.datac(\am_writing~q ),
	.datad(\wdata_burst_count[1]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~45_combout ),
	.cout());
defparam \p_main_fsm~45 .lut_mask = 16'hFFFE;
defparam \p_main_fsm~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~19 (
	.dataa(\state.s_idle~q ),
	.datab(\size_last[1]~q ),
	.datac(gnd),
	.datad(\rdata_bcount_eq_1~q ),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
defparam \Selector0~19 .lut_mask = 16'hEEFF;
defparam \Selector0~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~12 (
	.dataa(\Selector12~7_combout ),
	.datab(\p_main_fsm~45_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector53~12_combout ),
	.cout());
defparam \Selector53~12 .lut_mask = 16'hFEFF;
defparam \Selector53~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~13 (
	.dataa(\Selector42~11_combout ),
	.datab(\Selector12~4_combout ),
	.datac(\Selector53~11_combout ),
	.datad(\Selector53~12_combout ),
	.cin(gnd),
	.combout(\Selector53~13_combout ),
	.cout());
defparam \Selector53~13 .lut_mask = 16'hFFFE;
defparam \Selector53~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~14 (
	.dataa(\Selector12~9_combout ),
	.datab(\Selector53~10_combout ),
	.datac(\p_main_fsm~156_combout ),
	.datad(\Selector53~13_combout ),
	.cin(gnd),
	.combout(\Selector53~14_combout ),
	.cout());
defparam \Selector53~14 .lut_mask = 16'hFFFE;
defparam \Selector53~14 .sum_lutc_input = "datac";

dffeas didnt_write(
	.clk(clk),
	.d(\Selector53~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\didnt_write~q ),
	.prn(vcc));
defparam didnt_write.is_wysiwyg = "true";
defparam didnt_write.power_up = "low";

cycloneiii_lcell_comb \Selector4~4 (
	.dataa(\state.s_writing~q ),
	.datab(gnd),
	.datac(\write_req_this~q ),
	.datad(\didnt_write~q ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
defparam \Selector4~4 .lut_mask = 16'hAFFF;
defparam \Selector4~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state.s_wait_for_init_done~1 (
	.dataa(ctl_init_success),
	.datab(\state.s_wait_for_init_done~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state.s_wait_for_init_done~1_combout ),
	.cout());
defparam \state.s_wait_for_init_done~1 .lut_mask = 16'hEEEE;
defparam \state.s_wait_for_init_done~1 .sum_lutc_input = "datac";

dffeas \state.s_wait_for_init_done (
	.clk(clk),
	.d(\state.s_wait_for_init_done~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_wait_for_init_done~q ),
	.prn(vcc));
defparam \state.s_wait_for_init_done .is_wysiwyg = "true";
defparam \state.s_wait_for_init_done .power_up = "low";

cycloneiii_lcell_comb \Selector4~5 (
	.dataa(\Selector0~21_combout ),
	.datab(\Selector4~4_combout ),
	.datac(ctl_init_success),
	.datad(\state.s_wait_for_init_done~q ),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
defparam \Selector4~5 .lut_mask = 16'hFEFF;
defparam \Selector4~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~6 (
	.dataa(\state~331_combout ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
defparam \Selector4~6 .lut_mask = 16'hBFFF;
defparam \Selector4~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~7 (
	.dataa(\Selector4~3_combout ),
	.datab(\Selector4~5_combout ),
	.datac(\state.s_idle~q ),
	.datad(\Selector4~6_combout ),
	.cin(gnd),
	.combout(\Selector4~7_combout ),
	.cout());
defparam \Selector4~7 .lut_mask = 16'hFFFE;
defparam \Selector4~7 .sum_lutc_input = "datac";

dffeas \state.s_idle (
	.clk(clk),
	.d(\Selector4~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_idle~q ),
	.prn(vcc));
defparam \state.s_idle .is_wysiwyg = "true";
defparam \state.s_idle .power_up = "low";

cycloneiii_lcell_comb \Selector20~19 (
	.dataa(\size_last[1]~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\state.s_idle~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector20~19_combout ),
	.cout());
defparam \Selector20~19 .lut_mask = 16'hFBFF;
defparam \Selector20~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector39~0 (
	.dataa(\Selector5~6_combout ),
	.datab(\Selector20~19_combout ),
	.datac(\Selector20~2_combout ),
	.datad(\p_main_fsm~170_combout ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
defparam \Selector39~0 .lut_mask = 16'hFEFF;
defparam \Selector39~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector39~1 (
	.dataa(\new_req~q ),
	.datab(\read_req_this~q ),
	.datac(\write_req_this~q ),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\Selector39~1_combout ),
	.cout());
defparam \Selector39~1 .lut_mask = 16'hFEFF;
defparam \Selector39~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~7 (
	.dataa(\state.s_write~q ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\Selector5~7_combout ),
	.cout());
defparam \Selector5~7 .lut_mask = 16'hEFFF;
defparam \Selector5~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector39~2 (
	.dataa(\Selector26~0_combout ),
	.datab(\Selector39~0_combout ),
	.datac(\Selector39~1_combout ),
	.datad(\Selector5~7_combout ),
	.cin(gnd),
	.combout(\Selector39~2_combout ),
	.cout());
defparam \Selector39~2 .lut_mask = 16'hFFFD;
defparam \Selector39~2 .sum_lutc_input = "datac";

dffeas doing_act(
	.clk(clk),
	.d(\Selector39~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_act~q ),
	.prn(vcc));
defparam doing_act.is_wysiwyg = "true";
defparam doing_act.power_up = "low";

dffeas \trcd_pipe[0] (
	.clk(clk),
	.d(\doing_act~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trcd_pipe[0]~q ),
	.prn(vcc));
defparam \trcd_pipe[0] .is_wysiwyg = "true";
defparam \trcd_pipe[0] .power_up = "low";

dffeas finished_trcd(
	.clk(clk),
	.d(\trcd_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_trcd~q ),
	.prn(vcc));
defparam finished_trcd.is_wysiwyg = "true";
defparam finished_trcd.power_up = "low";

cycloneiii_lcell_comb \ba[1]~123 (
	.dataa(\state.s_activate~q ),
	.datab(\finished_trcd~q ),
	.datac(gnd),
	.datad(\doing_act~q ),
	.cin(gnd),
	.combout(\ba[1]~123_combout ),
	.cout());
defparam \ba[1]~123 .lut_mask = 16'hEEFF;
defparam \ba[1]~123 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~5 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\Selector20~19_combout ),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
defparam \Selector8~5 .lut_mask = 16'hFFFE;
defparam \Selector8~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~1 (
	.dataa(\p_main_fsm~39_combout ),
	.datab(\ba[1]~123_combout ),
	.datac(\p_main_fsm~63_combout ),
	.datad(\Selector8~5_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hFFFE;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~2 (
	.dataa(\Selector6~0_combout ),
	.datab(\read_req_this~q ),
	.datac(\Selector6~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hFEFE;
defparam \Selector6~2 .sum_lutc_input = "datac";

dffeas \state.s_read (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_read~q ),
	.prn(vcc));
defparam \state.s_read .is_wysiwyg = "true";
defparam \state.s_read .power_up = "low";

cycloneiii_lcell_comb \Selector20~4 (
	.dataa(\state.s_wait_for_init_done~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.s_refresh~q ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
defparam \Selector20~4 .lut_mask = 16'hAAFF;
defparam \Selector20~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~8 (
	.dataa(\state.s_precharge~q ),
	.datab(\state.s_read~q ),
	.datac(\state.s_holding~q ),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\Selector46~8_combout ),
	.cout());
defparam \Selector46~8 .lut_mask = 16'hFEFF;
defparam \Selector46~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \new_req~45 (
	.dataa(\rfsh_pending~q ),
	.datab(\in_buf|my_fifo|pipefull[0]~q ),
	.datac(\in_buf|my_fifo|pipe[0][28]~q ),
	.datad(\in_buf|my_fifo|pipe[0][27]~q ),
	.cin(gnd),
	.combout(\new_req~45_combout ),
	.cout());
defparam \new_req~45 .lut_mask = 16'hFFFE;
defparam \new_req~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \new_req~46 (
	.dataa(\accepted~q ),
	.datab(\accepted_r~q ),
	.datac(\size_last[1]~q ),
	.datad(\read_req_last~q ),
	.cin(gnd),
	.combout(\new_req~46_combout ),
	.cout());
defparam \new_req~46 .lut_mask = 16'hFFFE;
defparam \new_req~46 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \new_req~47 (
	.dataa(\new_req~q ),
	.datab(\new_req~45_combout ),
	.datac(\new_req~46_combout ),
	.datad(\read_req_last~2_combout ),
	.cin(gnd),
	.combout(\new_req~47_combout ),
	.cout());
defparam \new_req~47 .lut_mask = 16'hFEFF;
defparam \new_req~47 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~16 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector46~16_combout ),
	.cout());
defparam \Selector46~16 .lut_mask = 16'hFEFF;
defparam \Selector46~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~9 (
	.dataa(\state.s_write~q ),
	.datab(\read_req_this~q ),
	.datac(\p_main_fsm~105_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector46~9_combout ),
	.cout());
defparam \Selector46~9 .lut_mask = 16'hFFD8;
defparam \Selector46~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~10 (
	.dataa(\new_req~47_combout ),
	.datab(\Selector46~16_combout ),
	.datac(\state.s_write~q ),
	.datad(\Selector46~9_combout ),
	.cin(gnd),
	.combout(\Selector46~10_combout ),
	.cout());
defparam \Selector46~10 .lut_mask = 16'hFFFB;
defparam \Selector46~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~11 (
	.dataa(\process_13~0_combout ),
	.datab(\Selector46~8_combout ),
	.datac(\new_req~47_combout ),
	.datad(\Selector46~10_combout ),
	.cin(gnd),
	.combout(\Selector46~11_combout ),
	.cout());
defparam \Selector46~11 .lut_mask = 16'hFFFE;
defparam \Selector46~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_13~0 (
	.dataa(\accepted~q ),
	.datab(\in_buf|my_fifo|pipefull[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_13~0_combout ),
	.cout());
defparam \process_13~0 .lut_mask = 16'hEEEE;
defparam \process_13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~12 (
	.dataa(\Selector0~5_combout ),
	.datab(\Selector46~16_combout ),
	.datac(\ba[1]~122_combout ),
	.datad(\Selector43~0_combout ),
	.cin(gnd),
	.combout(\Selector46~12_combout ),
	.cout());
defparam \Selector46~12 .lut_mask = 16'hEFFF;
defparam \Selector46~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~13 (
	.dataa(\Selector46~7_combout ),
	.datab(\Selector46~11_combout ),
	.datac(\process_13~0_combout ),
	.datad(\Selector46~12_combout ),
	.cin(gnd),
	.combout(\Selector46~13_combout ),
	.cout());
defparam \Selector46~13 .lut_mask = 16'hFFFE;
defparam \Selector46~13 .sum_lutc_input = "datac";

dffeas new_req(
	.clk(clk),
	.d(\Selector46~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\new_req~q ),
	.prn(vcc));
defparam new_req.is_wysiwyg = "true";
defparam new_req.power_up = "low";

cycloneiii_lcell_comb \Selector11~1 (
	.dataa(\this_row_is_open~q ),
	.datab(\bank_is_open~q ),
	.datac(\new_req~q ),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
defparam \Selector11~1 .lut_mask = 16'hFEFF;
defparam \Selector11~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \new_req~49 (
	.dataa(\read_req_this~q ),
	.datab(\rdata_bcount_eq_0~q ),
	.datac(\finished_twtr~q ),
	.datad(\dqs_toggle_le_1~q ),
	.cin(gnd),
	.combout(\new_req~49_combout ),
	.cout());
defparam \new_req~49 .lut_mask = 16'hEFFF;
defparam \new_req~49 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~2 (
	.dataa(\ba[1]~123_combout ),
	.datab(\Selector37~2_combout ),
	.datac(\Selector11~1_combout ),
	.datad(\new_req~49_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
defparam \Selector11~2 .lut_mask = 16'hFFFE;
defparam \Selector11~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~20 (
	.dataa(\read_req_this~q ),
	.datab(\write_req_this~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~20_combout ),
	.cout());
defparam \p_main_fsm~20 .lut_mask = 16'hEEEE;
defparam \p_main_fsm~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~4 (
	.dataa(\new_req~q ),
	.datab(\state.s_write~q ),
	.datac(\p_main_fsm~20_combout ),
	.datad(\Selector44~15_combout ),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
defparam \Selector11~4 .lut_mask = 16'hFFFE;
defparam \Selector11~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~5 (
	.dataa(\Selector11~3_combout ),
	.datab(\Selector11~4_combout ),
	.datac(\Selector2~14_combout ),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
defparam \Selector11~5 .lut_mask = 16'hFEFF;
defparam \Selector11~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~6 (
	.dataa(\Selector11~0_combout ),
	.datab(\Selector11~2_combout ),
	.datac(\p_main_fsm~156_combout ),
	.datad(\Selector11~5_combout ),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
defparam \Selector11~6 .lut_mask = 16'hFFFE;
defparam \Selector11~6 .sum_lutc_input = "datac";

dffeas \state.s_reading (
	.clk(clk),
	.d(\Selector11~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_reading~q ),
	.prn(vcc));
defparam \state.s_reading .is_wysiwyg = "true";
defparam \state.s_reading .power_up = "low";

cycloneiii_lcell_comb \ba[1]~119 (
	.dataa(\a[5]~574_combout ),
	.datab(\cs_addr_to_term[0]~q ),
	.datac(gnd),
	.datad(\read_req_last~q ),
	.cin(gnd),
	.combout(\ba[1]~119_combout ),
	.cout());
defparam \ba[1]~119 .lut_mask = 16'hEEFF;
defparam \ba[1]~119 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~10 (
	.dataa(\p_main_fsm~156_combout ),
	.datab(\p_main_fsm~158_combout ),
	.datac(\ba[1]~118_combout ),
	.datad(\ba[1]~119_combout ),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
defparam \Selector0~10 .lut_mask = 16'hFFFE;
defparam \Selector0~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~11 (
	.dataa(\rdata_bcount_eq_1~q ),
	.datab(\didnt_term~q ),
	.datac(\new_req~q ),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
defparam \Selector0~11 .lut_mask = 16'hFFEF;
defparam \Selector0~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~12 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\rfsh_pending~q ),
	.datac(\state.s_reading~q ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
defparam \Selector0~12 .lut_mask = 16'hFFFB;
defparam \Selector0~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~17 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rfsh_pending~q ),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
defparam \Selector0~17 .lut_mask = 16'hAAFF;
defparam \Selector0~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~21 (
	.dataa(\state.s_refresh~q ),
	.datab(\finished_trfc~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
defparam \Selector0~21 .lut_mask = 16'hEEEE;
defparam \Selector0~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~22 (
	.dataa(\Selector0~20_combout ),
	.datab(\Selector0~21_combout ),
	.datac(\p_main_fsm~20_combout ),
	.datad(\new_req~q ),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
defparam \Selector0~22 .lut_mask = 16'hEFFF;
defparam \Selector0~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~23 (
	.dataa(\Selector0~16_combout ),
	.datab(\Selector0~17_combout ),
	.datac(\Selector0~22_combout ),
	.datad(\accepted~q ),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
defparam \Selector0~23 .lut_mask = 16'hFEFF;
defparam \Selector0~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~4 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][29]~q ),
	.datac(gnd),
	.datad(\rfsh_pending~q ),
	.cin(gnd),
	.combout(\Selector0~4_combout ),
	.cout());
defparam \Selector0~4 .lut_mask = 16'hEEFF;
defparam \Selector0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~25 (
	.dataa(\Selector0~24_combout ),
	.datab(\write_req_next~0_combout ),
	.datac(\Selector0~4_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
defparam \Selector0~25 .lut_mask = 16'hFFFE;
defparam \Selector0~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~26 (
	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector0~23_combout ),
	.datad(\Selector0~25_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
defparam \Selector0~26 .lut_mask = 16'hFFFE;
defparam \Selector0~26 .sum_lutc_input = "datac";

dffeas accepted(
	.clk(clk),
	.d(\Selector0~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\accepted~q ),
	.prn(vcc));
defparam accepted.is_wysiwyg = "true";
defparam accepted.power_up = "low";

dffeas read_req_this(
	.clk(clk),
	.d(\read_req_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\read_req_this~q ),
	.prn(vcc));
defparam read_req_this.is_wysiwyg = "true";
defparam read_req_this.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~157 (
	.dataa(\new_req~q ),
	.datab(\read_req_this~q ),
	.datac(\write_req_this~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~157_combout ),
	.cout());
defparam \p_main_fsm~157 .lut_mask = 16'hFEFE;
defparam \p_main_fsm~157 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~332 (
	.dataa(\p_main_fsm~156_combout ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\state~332_combout ),
	.cout());
defparam \state~332 .lut_mask = 16'hEFFF;
defparam \state~332 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \am_writing~24 (
	.dataa(\wdata_burst_count[0]~q ),
	.datab(gnd),
	.datac(\am_writing~q ),
	.datad(\wdata_burst_count[1]~q ),
	.cin(gnd),
	.combout(\am_writing~24_combout ),
	.cout());
defparam \am_writing~24 .lut_mask = 16'hAFFF;
defparam \am_writing~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~1 (
	.dataa(\Selector50~0_combout ),
	.datab(\state~332_combout ),
	.datac(\wdata_burst_count[1]~51_combout ),
	.datad(\am_writing~24_combout ),
	.cin(gnd),
	.combout(\Selector50~1_combout ),
	.cout());
defparam \Selector50~1 .lut_mask = 16'hBFFF;
defparam \Selector50~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~2 (
	.dataa(\state.s_write~q ),
	.datab(\p_main_fsm~105_combout ),
	.datac(\am_writing~24_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector50~2_combout ),
	.cout());
defparam \Selector50~2 .lut_mask = 16'hBFFF;
defparam \Selector50~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~3 (
	.dataa(\Selector0~19_combout ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\p_main_fsm~45_combout ),
	.datad(\am_writing~24_combout ),
	.cin(gnd),
	.combout(\Selector50~3_combout ),
	.cout());
defparam \Selector50~3 .lut_mask = 16'hBFFF;
defparam \Selector50~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~4 (
	.dataa(\p_main_fsm~166_combout ),
	.datab(\Selector50~2_combout ),
	.datac(\Selector50~3_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector50~4_combout ),
	.cout());
defparam \Selector50~4 .lut_mask = 16'hFEFF;
defparam \Selector50~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~6 (
	.dataa(\finished_trcd~q ),
	.datab(\Selector50~5_combout ),
	.datac(\read_req_this~q ),
	.datad(\doing_act~q ),
	.cin(gnd),
	.combout(\Selector50~6_combout ),
	.cout());
defparam \Selector50~6 .lut_mask = 16'hEFFF;
defparam \Selector50~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~7 (
	.dataa(\state.s_activate~q ),
	.datab(\Selector50~6_combout ),
	.datac(gnd),
	.datad(\am_writing~24_combout ),
	.cin(gnd),
	.combout(\Selector50~7_combout ),
	.cout());
defparam \Selector50~7 .lut_mask = 16'hEEFF;
defparam \Selector50~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~8 (
	.dataa(\Selector8~2_combout ),
	.datab(\Selector50~1_combout ),
	.datac(\Selector50~4_combout ),
	.datad(\Selector50~7_combout ),
	.cin(gnd),
	.combout(\Selector50~8_combout ),
	.cout());
defparam \Selector50~8 .lut_mask = 16'hFFFE;
defparam \Selector50~8 .sum_lutc_input = "datac";

dffeas am_writing(
	.clk(clk),
	.d(\Selector50~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\am_writing~q ),
	.prn(vcc));
defparam am_writing.is_wysiwyg = "true";
defparam am_writing.power_up = "low";

cycloneiii_lcell_comb \Selector3~4 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\am_writing~q ),
	.datac(\writing_in_proc~q ),
	.datad(\bank_man|Equal8~0_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
defparam \Selector3~4 .lut_mask = 16'hFFBF;
defparam \Selector3~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dqs_toggle_eq_0~1 (
	.dataa(\state.s_write~q ),
	.datab(\dqs_must_keep_toggling[2]~q ),
	.datac(\dqs_must_keep_toggling[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\dqs_toggle_eq_0~1_combout ),
	.cout());
defparam \dqs_toggle_eq_0~1 .lut_mask = 16'hFEFE;
defparam \dqs_toggle_eq_0~1 .sum_lutc_input = "datac";

dffeas dqs_toggle_eq_0(
	.clk(clk),
	.d(\dqs_toggle_eq_0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_toggle_eq_0~q ),
	.prn(vcc));
defparam dqs_toggle_eq_0.is_wysiwyg = "true";
defparam dqs_toggle_eq_0.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~162 (
	.dataa(\p_main_fsm~161_combout ),
	.datab(\g_timers:3:bank_timer|twr_pipe[2]~q ),
	.datac(\g_timers:1:bank_timer|twr_pipe[2]~q ),
	.datad(\g_timers:0:bank_timer|twr_pipe[2]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~162_combout ),
	.cout());
defparam \p_main_fsm~162 .lut_mask = 16'hBFFF;
defparam \p_main_fsm~162 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal19~0 (
	.dataa(\g_timers:1:bank_timer|finished_tras~q ),
	.datab(\g_timers:2:bank_timer|finished_tras~q ),
	.datac(\g_timers:0:bank_timer|finished_tras~q ),
	.datad(\g_timers:3:bank_timer|finished_tras~q ),
	.cin(gnd),
	.combout(\Equal19~0_combout ),
	.cout());
defparam \Equal19~0 .lut_mask = 16'hFFFE;
defparam \Equal19~0 .sum_lutc_input = "datac";

dffeas finished_tras_all(
	.clk(clk),
	.d(\Equal19~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_tras_all~q ),
	.prn(vcc));
defparam finished_tras_all.is_wysiwyg = "true";
defparam finished_tras_all.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~163 (
	.dataa(\p_main_fsm~160_combout ),
	.datab(\dqs_toggle_eq_0~q ),
	.datac(\p_main_fsm~162_combout ),
	.datad(\finished_tras_all~q ),
	.cin(gnd),
	.combout(\p_main_fsm~163_combout ),
	.cout());
defparam \p_main_fsm~163 .lut_mask = 16'hEFFF;
defparam \p_main_fsm~163 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector23~3 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\bank_man|Equal8~0_combout ),
	.datad(\p_main_fsm~163_combout ),
	.cin(gnd),
	.combout(\Selector23~3_combout ),
	.cout());
defparam \Selector23~3 .lut_mask = 16'hEFFF;
defparam \Selector23~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector21~0 (
	.dataa(\refresh_in_progress~q ),
	.datab(\Selector23~3_combout ),
	.datac(\state.s_refresh~q ),
	.datad(\finished_trfc~q ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
defparam \Selector21~0 .lut_mask = 16'hACFF;
defparam \Selector21~0 .sum_lutc_input = "datac";

dffeas refresh_in_progress(
	.clk(clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_in_progress~q ),
	.prn(vcc));
defparam refresh_in_progress.is_wysiwyg = "true";
defparam refresh_in_progress.power_up = "low";

cycloneiii_lcell_comb \p_main_fsm~57 (
	.dataa(\rfsh_pending~q ),
	.datab(\refresh_in_progress~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~57_combout ),
	.cout());
defparam \p_main_fsm~57 .lut_mask = 16'hEEEE;
defparam \p_main_fsm~57 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(\bank_addr_this[1]~q ),
	.datab(\g_timers:1:bank_timer|finished_twr~combout ),
	.datac(\bank_addr_this[0]~q ),
	.datad(\g_timers:0:bank_timer|finished_twr~combout ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~1 (
	.dataa(\g_timers:2:bank_timer|finished_twr~combout ),
	.datab(\bank_addr_this[1]~q ),
	.datac(\Mux2~0_combout ),
	.datad(\g_timers:3:bank_timer|finished_twr~combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~7 (
	.dataa(\am_writing~q ),
	.datab(\am_reading~q ),
	.datac(\finished_tras_all~q ),
	.datad(\Mux2~1_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
defparam \Selector2~7 .lut_mask = 16'hFFF7;
defparam \Selector2~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~8 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\p_main_fsm~163_combout ),
	.datad(\Selector2~7_combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
defparam \Selector2~8 .lut_mask = 16'hBF8F;
defparam \Selector2~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~13 (
	.dataa(\state.s_holding~q ),
	.datab(\didnt_act~q ),
	.datac(\didnt_pch~q ),
	.datad(\p_main_fsm~165_combout ),
	.cin(gnd),
	.combout(\Selector2~13_combout ),
	.cout());
defparam \Selector2~13 .lut_mask = 16'hFBFF;
defparam \Selector2~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~9 (
	.dataa(\state~328_combout ),
	.datab(\Selector20~2_combout ),
	.datac(\finished_tras~q ),
	.datad(\finished_tras_last~q ),
	.cin(gnd),
	.combout(\Selector2~9_combout ),
	.cout());
defparam \Selector2~9 .lut_mask = 16'hFFFE;
defparam \Selector2~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~10 (
	.dataa(\p_main_fsm~157_combout ),
	.datab(\Mux2~1_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\Selector2~9_combout ),
	.cin(gnd),
	.combout(\Selector2~10_combout ),
	.cout());
defparam \Selector2~10 .lut_mask = 16'hFFFE;
defparam \Selector2~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~11 (
	.dataa(\Selector2~6_combout ),
	.datab(\Selector2~8_combout ),
	.datac(\Selector2~13_combout ),
	.datad(\Selector2~10_combout ),
	.cin(gnd),
	.combout(\Selector2~11_combout ),
	.cout());
defparam \Selector2~11 .lut_mask = 16'hFFFE;
defparam \Selector2~11 .sum_lutc_input = "datac";

dffeas doing_pch(
	.clk(clk),
	.d(\Selector2~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_pch~q ),
	.prn(vcc));
defparam doing_pch.is_wysiwyg = "true";
defparam doing_pch.power_up = "low";

dffeas \trp_pipe[0] (
	.clk(clk),
	.d(\doing_pch~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trp_pipe[0]~q ),
	.prn(vcc));
defparam \trp_pipe[0] .is_wysiwyg = "true";
defparam \trp_pipe[0] .power_up = "low";

dffeas finished_trp(
	.clk(clk),
	.d(\trp_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_trp~q ),
	.prn(vcc));
defparam finished_trp.is_wysiwyg = "true";
defparam finished_trp.power_up = "low";

cycloneiii_lcell_comb \Selector5~2 (
	.dataa(\state.s_precharge~q ),
	.datab(\finished_trp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hEEEE;
defparam \Selector5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~2 (
	.dataa(\Selector23~2_combout ),
	.datab(\Selector3~4_combout ),
	.datac(\p_main_fsm~57_combout ),
	.datad(\Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hFFFE;
defparam \Selector3~2 .sum_lutc_input = "datac";

dffeas doing_rfsh(
	.clk(clk),
	.d(\Selector3~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_rfsh~q ),
	.prn(vcc));
defparam doing_rfsh.is_wysiwyg = "true";
defparam doing_rfsh.power_up = "low";

dffeas \trfc_pipe[0] (
	.clk(clk),
	.d(\doing_rfsh~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[0]~q ),
	.prn(vcc));
defparam \trfc_pipe[0] .is_wysiwyg = "true";
defparam \trfc_pipe[0] .power_up = "low";

dffeas \trfc_pipe[1] (
	.clk(clk),
	.d(\trfc_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[1]~q ),
	.prn(vcc));
defparam \trfc_pipe[1] .is_wysiwyg = "true";
defparam \trfc_pipe[1] .power_up = "low";

dffeas \trfc_pipe[2] (
	.clk(clk),
	.d(\trfc_pipe[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[2]~q ),
	.prn(vcc));
defparam \trfc_pipe[2] .is_wysiwyg = "true";
defparam \trfc_pipe[2] .power_up = "low";

dffeas \trfc_pipe[3] (
	.clk(clk),
	.d(\trfc_pipe[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[3]~q ),
	.prn(vcc));
defparam \trfc_pipe[3] .is_wysiwyg = "true";
defparam \trfc_pipe[3] .power_up = "low";

dffeas \trfc_pipe[4] (
	.clk(clk),
	.d(\trfc_pipe[3]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[4]~q ),
	.prn(vcc));
defparam \trfc_pipe[4] .is_wysiwyg = "true";
defparam \trfc_pipe[4] .power_up = "low";

dffeas \trfc_pipe[5] (
	.clk(clk),
	.d(\trfc_pipe[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[5]~q ),
	.prn(vcc));
defparam \trfc_pipe[5] .is_wysiwyg = "true";
defparam \trfc_pipe[5] .power_up = "low";

dffeas \trfc_pipe[6] (
	.clk(clk),
	.d(\trfc_pipe[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[6]~q ),
	.prn(vcc));
defparam \trfc_pipe[6] .is_wysiwyg = "true";
defparam \trfc_pipe[6] .power_up = "low";

dffeas \trfc_pipe[7] (
	.clk(clk),
	.d(\trfc_pipe[6]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trfc_pipe[7]~q ),
	.prn(vcc));
defparam \trfc_pipe[7] .is_wysiwyg = "true";
defparam \trfc_pipe[7] .power_up = "low";

dffeas finished_trfc(
	.clk(clk),
	.d(\trfc_pipe[7]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_trfc~q ),
	.prn(vcc));
defparam finished_trfc.is_wysiwyg = "true";
defparam finished_trfc.power_up = "low";

cycloneiii_lcell_comb \Selector3~3 (
	.dataa(\state.s_refresh~q ),
	.datab(gnd),
	.datac(\finished_trfc~q ),
	.datad(\Selector3~2_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'hFFAF;
defparam \Selector3~3 .sum_lutc_input = "datac";

dffeas \state.s_refresh (
	.clk(clk),
	.d(\Selector3~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_refresh~q ),
	.prn(vcc));
defparam \state.s_refresh .is_wysiwyg = "true";
defparam \state.s_refresh .power_up = "low";

cycloneiii_lcell_comb \Selector2~12 (
	.dataa(\state.s_precharge~q ),
	.datab(gnd),
	.datac(\finished_trp~q ),
	.datad(\Selector2~11_combout ),
	.cin(gnd),
	.combout(\Selector2~12_combout ),
	.cout());
defparam \Selector2~12 .lut_mask = 16'hFFAF;
defparam \Selector2~12 .sum_lutc_input = "datac";

dffeas \state.s_precharge (
	.clk(clk),
	.d(\Selector2~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_precharge~q ),
	.prn(vcc));
defparam \state.s_precharge .is_wysiwyg = "true";
defparam \state.s_precharge .power_up = "low";

cycloneiii_lcell_comb \ba[1]~116 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_precharge~q ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\ba[1]~116_combout ),
	.cout());
defparam \ba[1]~116 .lut_mask = 16'h0FFF;
defparam \ba[1]~116 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector15~0 (
	.dataa(\rfsh_done~q ),
	.datab(\state.s_refresh~q ),
	.datac(\ba[1]~116_combout ),
	.datad(\Selector3~2_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hFFBF;
defparam \Selector15~0 .sum_lutc_input = "datac";

dffeas rfsh_done(
	.clk(clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rfsh_done~q ),
	.prn(vcc));
defparam rfsh_done.is_wysiwyg = "true";
defparam rfsh_done.power_up = "low";

cycloneiii_lcell_comb \rdata_valid_pipe~2 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_read~q ),
	.datac(gnd),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\rdata_valid_pipe~2_combout ),
	.cout());
defparam \rdata_valid_pipe~2 .lut_mask = 16'hEEFF;
defparam \rdata_valid_pipe~2 .sum_lutc_input = "datac";

dffeas \rdata_valid_pipe[2] (
	.clk(clk),
	.d(\rdata_valid_pipe~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_valid_pipe[2]~q ),
	.prn(vcc));
defparam \rdata_valid_pipe[2] .is_wysiwyg = "true";
defparam \rdata_valid_pipe[2] .power_up = "low";

cycloneiii_lcell_comb \a[5]~576 (
	.dataa(\size_last[1]~q ),
	.datab(gnd),
	.datac(\rdata_bcount_eq_1~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\a[5]~576_combout ),
	.cout());
defparam \a[5]~576 .lut_mask = 16'hAFFF;
defparam \a[5]~576 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \new_req~48 (
	.dataa(\p_main_fsm~45_combout ),
	.datab(gnd),
	.datac(\read_req_this~q ),
	.datad(\p_main_fsm~39_combout ),
	.cin(gnd),
	.combout(\new_req~48_combout ),
	.cout());
defparam \new_req~48 .lut_mask = 16'hA0AF;
defparam \new_req~48 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~2 (
	.dataa(\Selector17~1_combout ),
	.datab(\p_main_fsm~156_combout ),
	.datac(\a[5]~576_combout ),
	.datad(\new_req~48_combout ),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
defparam \Selector17~2 .lut_mask = 16'hFFFE;
defparam \Selector17~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \cs_n~61 (
	.dataa(\am_reading~q ),
	.datab(\finished_tras_all~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cs_n~61_combout ),
	.cout());
defparam \cs_n~61 .lut_mask = 16'hBBBB;
defparam \cs_n~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \cs_n~62 (
	.dataa(\state~328_combout ),
	.datab(\am_writing~q ),
	.datac(\Mux2~1_combout ),
	.datad(\cs_n~61_combout ),
	.cin(gnd),
	.combout(\cs_n~62_combout ),
	.cout());
defparam \cs_n~62 .lut_mask = 16'hFFEF;
defparam \cs_n~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~3 (
	.dataa(\state~331_combout ),
	.datab(\Selector17~2_combout ),
	.datac(\a[5]~576_combout ),
	.datad(\cs_n~62_combout ),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
defparam \Selector17~3 .lut_mask = 16'hFFFE;
defparam \Selector17~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~6 (
	.dataa(\Selector17~4_combout ),
	.datab(\Selector17~5_combout ),
	.datac(\state.s_holding~q ),
	.datad(\Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
defparam \Selector17~6 .lut_mask = 16'hEFFF;
defparam \Selector17~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector0~18 (
	.dataa(\size_last[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\size_last[1]~q ),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
defparam \Selector0~18 .lut_mask = 16'hAAFF;
defparam \Selector0~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~333 (
	.dataa(\size_last[1]~q ),
	.datab(\new_req~q ),
	.datac(\read_req_this~q ),
	.datad(\write_req_this~q ),
	.cin(gnd),
	.combout(\state~333_combout ),
	.cout());
defparam \state~333 .lut_mask = 16'hFFFE;
defparam \state~333 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~8 (
	.dataa(\Selector17~7_combout ),
	.datab(\Selector0~18_combout ),
	.datac(\state~333_combout ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\Selector17~8_combout ),
	.cout());
defparam \Selector17~8 .lut_mask = 16'hBFFF;
defparam \Selector17~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~169 (
	.dataa(\read_req_this~q ),
	.datab(\didnt_read~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\p_main_fsm~169_combout ),
	.cout());
defparam \p_main_fsm~169 .lut_mask = 16'hEEEE;
defparam \p_main_fsm~169 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~9 (
	.dataa(\didnt_term~q ),
	.datab(\read_req_last~q ),
	.datac(\cs_addr_to_term[0]~q ),
	.datad(\state.s_reading~q ),
	.cin(gnd),
	.combout(\Selector17~9_combout ),
	.cout());
defparam \Selector17~9 .lut_mask = 16'hEFFF;
defparam \Selector17~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~10 (
	.dataa(\didnt_term~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\a[5]~574_combout ),
	.datad(\Selector17~9_combout ),
	.cin(gnd),
	.combout(\Selector17~10_combout ),
	.cout());
defparam \Selector17~10 .lut_mask = 16'hBF1F;
defparam \Selector17~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~11 (
	.dataa(\didnt_term~q ),
	.datab(\p_main_fsm~169_combout ),
	.datac(\p_main_fsm~158_combout ),
	.datad(\Selector17~10_combout ),
	.cin(gnd),
	.combout(\Selector17~11_combout ),
	.cout());
defparam \Selector17~11 .lut_mask = 16'hF7B3;
defparam \Selector17~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~12 (
	.dataa(\size_last[1]~q ),
	.datab(\state.s_reading~q ),
	.datac(\Selector17~11_combout ),
	.datad(\Selector17~8_combout ),
	.cin(gnd),
	.combout(\Selector17~12_combout ),
	.cout());
defparam \Selector17~12 .lut_mask = 16'hFFFB;
defparam \Selector17~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~13 (
	.dataa(\cs_n~63_combout ),
	.datab(\cs_n~64_combout ),
	.datac(\Selector17~8_combout ),
	.datad(\Selector17~12_combout ),
	.cin(gnd),
	.combout(\Selector17~13_combout ),
	.cout());
defparam \Selector17~13 .lut_mask = 16'hFFFE;
defparam \Selector17~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~15 (
	.dataa(\bank_is_open~q ),
	.datab(\read_req_this~q ),
	.datac(\p_main_fsm~105_combout ),
	.datad(\this_row_is_open~q ),
	.cin(gnd),
	.combout(\Selector17~15_combout ),
	.cout());
defparam \Selector17~15 .lut_mask = 16'hFEFF;
defparam \Selector17~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~3 (
	.dataa(\state.s_write~q ),
	.datab(\p_main_fsm~157_combout ),
	.datac(gnd),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector42~3_combout ),
	.cout());
defparam \Selector42~3 .lut_mask = 16'hEEFF;
defparam \Selector42~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~16 (
	.dataa(\Selector17~14_combout ),
	.datab(\Selector17~15_combout ),
	.datac(\Selector42~3_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(\Selector17~16_combout ),
	.cout());
defparam \Selector17~16 .lut_mask = 16'hEFFF;
defparam \Selector17~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~17 (
	.dataa(\Selector17~3_combout ),
	.datab(\Selector17~6_combout ),
	.datac(\Selector17~13_combout ),
	.datad(\Selector17~16_combout ),
	.cin(gnd),
	.combout(\Selector17~17_combout ),
	.cout());
defparam \Selector17~17 .lut_mask = 16'h7FFF;
defparam \Selector17~17 .sum_lutc_input = "datac";

dffeas \row_addr_this[0] (
	.clk(clk),
	.d(\row_addr_next[0]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[0]~q ),
	.prn(vcc));
defparam \row_addr_this[0] .is_wysiwyg = "true";
defparam \row_addr_this[0] .power_up = "low";

cycloneiii_lcell_comb \a[0]~582 (
	.dataa(\finished_trp~q ),
	.datab(\state.s_precharge~q ),
	.datac(\bank_is_open~q ),
	.datad(\Selector37~2_combout ),
	.cin(gnd),
	.combout(\a[0]~582_combout ),
	.cout());
defparam \a[0]~582 .lut_mask = 16'h8BFF;
defparam \a[0]~582 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~583 (
	.dataa(\a[0]~581_combout ),
	.datab(\state.s_write~q ),
	.datac(\a[0]~582_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\a[0]~583_combout ),
	.cout());
defparam \a[0]~583 .lut_mask = 16'hFEFF;
defparam \a[0]~583 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~584 (
	.dataa(\state.s_precharge~q ),
	.datab(\rfsh_pending~q ),
	.datac(\refresh_in_progress~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[5]~584_combout ),
	.cout());
defparam \a[5]~584 .lut_mask = 16'hFEFE;
defparam \a[5]~584 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~585 (
	.dataa(\p_main_fsm~157_combout ),
	.datab(gnd),
	.datac(\state.s_idle~q ),
	.datad(\a[5]~584_combout ),
	.cin(gnd),
	.combout(\a[0]~585_combout ),
	.cout());
defparam \a[0]~585 .lut_mask = 16'hAFFF;
defparam \a[0]~585 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~586 (
	.dataa(\state.s_precharge~q ),
	.datab(\state.s_idle~q ),
	.datac(\state.s_write~q ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\a[0]~586_combout ),
	.cout());
defparam \a[0]~586 .lut_mask = 16'h7FFF;
defparam \a[0]~586 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~587 (
	.dataa(\state.s_holding~q ),
	.datab(\a[0]~583_combout ),
	.datac(\a[0]~585_combout ),
	.datad(\a[0]~586_combout ),
	.cin(gnd),
	.combout(\a[0]~587_combout ),
	.cout());
defparam \a[0]~587 .lut_mask = 16'hFFFE;
defparam \a[0]~587 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~5 (
	.dataa(\state.s_idle~q ),
	.datab(\p_main_fsm~19_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\bank_is_open~q ),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
defparam \Selector20~5 .lut_mask = 16'hEFFF;
defparam \Selector20~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~588 (
	.dataa(\Selector5~6_combout ),
	.datab(\size_last[1]~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\a[0]~588_combout ),
	.cout());
defparam \a[0]~588 .lut_mask = 16'hFAFC;
defparam \a[0]~588 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~589 (
	.dataa(\a[0]~578_combout ),
	.datab(\a[0]~587_combout ),
	.datac(\Selector20~5_combout ),
	.datad(\a[0]~588_combout ),
	.cin(gnd),
	.combout(\a[0]~589_combout ),
	.cout());
defparam \a[0]~589 .lut_mask = 16'hFFFE;
defparam \a[0]~589 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~155 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(gnd),
	.datac(\am_writing~q ),
	.datad(\writing_in_proc~q ),
	.cin(gnd),
	.combout(\p_main_fsm~155_combout ),
	.cout());
defparam \p_main_fsm~155 .lut_mask = 16'hAFFF;
defparam \p_main_fsm~155 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[0]~590 (
	.dataa(\state.s_holding~q ),
	.datab(\changing_cs_pause~q ),
	.datac(\p_main_fsm~155_combout ),
	.datad(\didnt_act~q ),
	.cin(gnd),
	.combout(\a[0]~590_combout ),
	.cout());
defparam \a[0]~590 .lut_mask = 16'hEFFF;
defparam \a[0]~590 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector36~0 (
	.dataa(\row_addr_this[0]~q ),
	.datab(\a[0]~589_combout ),
	.datac(gnd),
	.datad(\a[0]~590_combout ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hEEFF;
defparam \Selector36~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[0]~0 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[0]~0_combout ),
	.cout());
defparam \col_addr_next[0]~0 .lut_mask = 16'hEEEE;
defparam \col_addr_next[0]~0 .sum_lutc_input = "datac";

dffeas \col_addr_this[0] (
	.clk(clk),
	.d(\col_addr_next[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[0]~q ),
	.prn(vcc));
defparam \col_addr_this[0] .is_wysiwyg = "true";
defparam \col_addr_this[0] .power_up = "low";

cycloneiii_lcell_comb \row_addr_next[1]~1 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[1]~1_combout ),
	.cout());
defparam \row_addr_next[1]~1 .lut_mask = 16'hEEEE;
defparam \row_addr_next[1]~1 .sum_lutc_input = "datac";

dffeas \row_addr_this[1] (
	.clk(clk),
	.d(\row_addr_next[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[1]~q ),
	.prn(vcc));
defparam \row_addr_this[1] .is_wysiwyg = "true";
defparam \row_addr_this[1] .power_up = "low";

cycloneiii_lcell_comb \a[5]~594 (
	.dataa(\state.s_activate~q ),
	.datab(\p_main_fsm~63_combout ),
	.datac(\Selector50~5_combout ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\a[5]~594_combout ),
	.cout());
defparam \a[5]~594 .lut_mask = 16'hFAFC;
defparam \a[5]~594 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~595 (
	.dataa(\ba[1]~117_combout ),
	.datab(\wdata_burst_count[1]~53_combout ),
	.datac(\a[5]~594_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\a[5]~595_combout ),
	.cout());
defparam \a[5]~595 .lut_mask = 16'hFEFF;
defparam \a[5]~595 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~597 (
	.dataa(\state.s_idle~q ),
	.datab(\bank_is_open~q ),
	.datac(\size_last[1]~q ),
	.datad(\rdata_bcount_eq_1~q ),
	.cin(gnd),
	.combout(\a[5]~597_combout ),
	.cout());
defparam \a[5]~597 .lut_mask = 16'hFEFF;
defparam \a[5]~597 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~598 (
	.dataa(\a[5]~596_combout ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\a[5]~597_combout ),
	.cin(gnd),
	.combout(\a[5]~598_combout ),
	.cout());
defparam \a[5]~598 .lut_mask = 16'hFFDF;
defparam \a[5]~598 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~127 (
	.dataa(\state.s_write~q ),
	.datab(\this_row_is_open~q ),
	.datac(\bank_is_open~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ba[1]~127_combout ),
	.cout());
defparam \ba[1]~127 .lut_mask = 16'h7F7F;
defparam \ba[1]~127 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~128 (
	.dataa(\p_main_fsm~154_combout ),
	.datab(\state.s_writing~q ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\ba[1]~127_combout ),
	.cin(gnd),
	.combout(\ba[1]~128_combout ),
	.cout());
defparam \ba[1]~128 .lut_mask = 16'hFFBF;
defparam \ba[1]~128 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdata_burst_count[1]~69 (
	.dataa(\read_req_this~q ),
	.datab(\state.s_writing~q ),
	.datac(\write_req_this~q ),
	.datad(\didnt_write~q ),
	.cin(gnd),
	.combout(\wdata_burst_count[1]~69_combout ),
	.cout());
defparam \wdata_burst_count[1]~69 .lut_mask = 16'h8BFF;
defparam \wdata_burst_count[1]~69 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~599 (
	.dataa(\ba[1]~123_combout ),
	.datab(\a[5]~598_combout ),
	.datac(\ba[1]~128_combout ),
	.datad(\wdata_burst_count[1]~69_combout ),
	.cin(gnd),
	.combout(\a[5]~599_combout ),
	.cout());
defparam \a[5]~599 .lut_mask = 16'hEFFF;
defparam \a[5]~599 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~600 (
	.dataa(\a[5]~593_combout ),
	.datab(\a[5]~595_combout ),
	.datac(\a[5]~599_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[5]~600_combout ),
	.cout());
defparam \a[5]~600 .lut_mask = 16'hFEFE;
defparam \a[5]~600 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~605 (
	.dataa(\a[5]~576_combout ),
	.datab(\Selector39~1_combout ),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\state.s_precharge~q ),
	.cin(gnd),
	.combout(\a[5]~605_combout ),
	.cout());
defparam \a[5]~605 .lut_mask = 16'hFFFE;
defparam \a[5]~605 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~575 (
	.dataa(\p_main_fsm~157_combout ),
	.datab(\size_last[1]~q ),
	.datac(\rdata_bcount_eq_1~q ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\a[5]~575_combout ),
	.cout());
defparam \a[5]~575 .lut_mask = 16'hEFFF;
defparam \a[5]~575 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~606 (
	.dataa(\a[5]~596_combout ),
	.datab(\bank_is_open~q ),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\a[5]~575_combout ),
	.cin(gnd),
	.combout(\a[5]~606_combout ),
	.cout());
defparam \a[5]~606 .lut_mask = 16'hF7D5;
defparam \a[5]~606 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~607 (
	.dataa(\am_writing~q ),
	.datab(\state.s_idle~q ),
	.datac(\a[5]~605_combout ),
	.datad(\a[5]~606_combout ),
	.cin(gnd),
	.combout(\a[5]~607_combout ),
	.cout());
defparam \a[5]~607 .lut_mask = 16'hFEFF;
defparam \a[5]~607 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~596 (
	.dataa(\state.s_activate~q ),
	.datab(\doing_act~q ),
	.datac(\finished_trcd~q ),
	.datad(\this_row_is_open~q ),
	.cin(gnd),
	.combout(\a[5]~596_combout ),
	.cout());
defparam \a[5]~596 .lut_mask = 16'h8DFF;
defparam \a[5]~596 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~609 (
	.dataa(\a[0]~590_combout ),
	.datab(\state.s_activate~q ),
	.datac(\a[5]~596_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\a[5]~609_combout ),
	.cout());
defparam \a[5]~609 .lut_mask = 16'hFEFE;
defparam \a[5]~609 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~610 (
	.dataa(\a[5]~608_combout ),
	.datab(\a[5]~609_combout ),
	.datac(\wdata_burst_count[1]~69_combout ),
	.datad(\ba[1]~128_combout ),
	.cin(gnd),
	.combout(\a[5]~610_combout ),
	.cout());
defparam \a[5]~610 .lut_mask = 16'hFEFF;
defparam \a[5]~610 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~612 (
	.dataa(\Selector37~2_combout ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\state.s_write~q ),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\a[5]~612_combout ),
	.cout());
defparam \a[5]~612 .lut_mask = 16'hFEFF;
defparam \a[5]~612 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~126 (
	.dataa(\size_last[1]~q ),
	.datab(\write_req_this~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ba[1]~126_combout ),
	.cout());
defparam \ba[1]~126 .lut_mask = 16'hEEEE;
defparam \ba[1]~126 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~592 (
	.dataa(\p_main_fsm~168_combout ),
	.datab(\ba[1]~126_combout ),
	.datac(\state.s_reading~q ),
	.datad(\a[5]~574_combout ),
	.cin(gnd),
	.combout(\a[5]~592_combout ),
	.cout());
defparam \a[5]~592 .lut_mask = 16'hACFF;
defparam \a[5]~592 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~591 (
	.dataa(\size_last[1]~q ),
	.datab(\p_main_fsm~156_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\state.s_read~q ),
	.cin(gnd),
	.combout(\a[5]~591_combout ),
	.cout());
defparam \a[5]~591 .lut_mask = 16'hFFFE;
defparam \a[5]~591 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~613 (
	.dataa(\a[5]~611_combout ),
	.datab(\a[5]~612_combout ),
	.datac(\a[5]~592_combout ),
	.datad(\a[5]~591_combout ),
	.cin(gnd),
	.combout(\a[5]~613_combout ),
	.cout());
defparam \a[5]~613 .lut_mask = 16'hFFFE;
defparam \a[5]~613 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \a[5]~614 (
	.dataa(\a[5]~604_combout ),
	.datab(\a[5]~607_combout ),
	.datac(\a[5]~610_combout ),
	.datad(\a[5]~613_combout ),
	.cin(gnd),
	.combout(\a[5]~614_combout ),
	.cout());
defparam \a[5]~614 .lut_mask = 16'hFFFE;
defparam \a[5]~614 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector35~0 (
	.dataa(\col_addr_this[0]~q ),
	.datab(\row_addr_this[1]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector35~0_combout ),
	.cout());
defparam \Selector35~0 .lut_mask = 16'hACFF;
defparam \Selector35~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[1]~1 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[1]~1_combout ),
	.cout());
defparam \col_addr_next[1]~1 .lut_mask = 16'hEEEE;
defparam \col_addr_next[1]~1 .sum_lutc_input = "datac";

dffeas \col_addr_this[1] (
	.clk(clk),
	.d(\col_addr_next[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[1]~q ),
	.prn(vcc));
defparam \col_addr_this[1] .is_wysiwyg = "true";
defparam \col_addr_this[1] .power_up = "low";

dffeas \row_addr_this[2] (
	.clk(clk),
	.d(\row_addr_next[2]~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[2]~q ),
	.prn(vcc));
defparam \row_addr_this[2] .is_wysiwyg = "true";
defparam \row_addr_this[2] .power_up = "low";

cycloneiii_lcell_comb \Selector34~0 (
	.dataa(\col_addr_this[1]~q ),
	.datab(\row_addr_this[2]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector34~0_combout ),
	.cout());
defparam \Selector34~0 .lut_mask = 16'hACFF;
defparam \Selector34~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[2]~2 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[2]~2_combout ),
	.cout());
defparam \col_addr_next[2]~2 .lut_mask = 16'hEEEE;
defparam \col_addr_next[2]~2 .sum_lutc_input = "datac";

dffeas \col_addr_this[2] (
	.clk(clk),
	.d(\col_addr_next[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[2]~q ),
	.prn(vcc));
defparam \col_addr_this[2] .is_wysiwyg = "true";
defparam \col_addr_this[2] .power_up = "low";

dffeas \row_addr_this[3] (
	.clk(clk),
	.d(\row_addr_next[3]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[3]~q ),
	.prn(vcc));
defparam \row_addr_this[3] .is_wysiwyg = "true";
defparam \row_addr_this[3] .power_up = "low";

cycloneiii_lcell_comb \Selector33~0 (
	.dataa(\col_addr_this[2]~q ),
	.datab(\row_addr_this[3]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'hACFF;
defparam \Selector33~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[3]~3 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[3]~3_combout ),
	.cout());
defparam \col_addr_next[3]~3 .lut_mask = 16'hEEEE;
defparam \col_addr_next[3]~3 .sum_lutc_input = "datac";

dffeas \col_addr_this[3] (
	.clk(clk),
	.d(\col_addr_next[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[3]~q ),
	.prn(vcc));
defparam \col_addr_this[3] .is_wysiwyg = "true";
defparam \col_addr_this[3] .power_up = "low";

cycloneiii_lcell_comb \row_addr_next[4]~2 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[4]~2_combout ),
	.cout());
defparam \row_addr_next[4]~2 .lut_mask = 16'hEEEE;
defparam \row_addr_next[4]~2 .sum_lutc_input = "datac";

dffeas \row_addr_this[4] (
	.clk(clk),
	.d(\row_addr_next[4]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[4]~q ),
	.prn(vcc));
defparam \row_addr_this[4] .is_wysiwyg = "true";
defparam \row_addr_this[4] .power_up = "low";

cycloneiii_lcell_comb \Selector32~0 (
	.dataa(\col_addr_this[3]~q ),
	.datab(\row_addr_this[4]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'hACFF;
defparam \Selector32~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[4]~4 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[4]~4_combout ),
	.cout());
defparam \col_addr_next[4]~4 .lut_mask = 16'hEEEE;
defparam \col_addr_next[4]~4 .sum_lutc_input = "datac";

dffeas \col_addr_this[4] (
	.clk(clk),
	.d(\col_addr_next[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[4]~q ),
	.prn(vcc));
defparam \col_addr_this[4] .is_wysiwyg = "true";
defparam \col_addr_this[4] .power_up = "low";

dffeas \row_addr_this[5] (
	.clk(clk),
	.d(\row_addr_next[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[5]~q ),
	.prn(vcc));
defparam \row_addr_this[5] .is_wysiwyg = "true";
defparam \row_addr_this[5] .power_up = "low";

cycloneiii_lcell_comb \Selector31~0 (
	.dataa(\col_addr_this[4]~q ),
	.datab(\row_addr_this[5]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
defparam \Selector31~0 .lut_mask = 16'hACFF;
defparam \Selector31~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[5]~5 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[5]~5_combout ),
	.cout());
defparam \col_addr_next[5]~5 .lut_mask = 16'hEEEE;
defparam \col_addr_next[5]~5 .sum_lutc_input = "datac";

dffeas \col_addr_this[5] (
	.clk(clk),
	.d(\col_addr_next[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[5]~q ),
	.prn(vcc));
defparam \col_addr_this[5] .is_wysiwyg = "true";
defparam \col_addr_this[5] .power_up = "low";

cycloneiii_lcell_comb \row_addr_next[6]~7 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[6]~7_combout ),
	.cout());
defparam \row_addr_next[6]~7 .lut_mask = 16'hEEEE;
defparam \row_addr_next[6]~7 .sum_lutc_input = "datac";

dffeas \row_addr_this[6] (
	.clk(clk),
	.d(\row_addr_next[6]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[6]~q ),
	.prn(vcc));
defparam \row_addr_this[6] .is_wysiwyg = "true";
defparam \row_addr_this[6] .power_up = "low";

cycloneiii_lcell_comb \Selector30~0 (
	.dataa(\col_addr_this[5]~q ),
	.datab(\row_addr_this[6]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
defparam \Selector30~0 .lut_mask = 16'hACFF;
defparam \Selector30~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[6]~6 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[6]~6_combout ),
	.cout());
defparam \col_addr_next[6]~6 .lut_mask = 16'hEEEE;
defparam \col_addr_next[6]~6 .sum_lutc_input = "datac";

dffeas \col_addr_this[6] (
	.clk(clk),
	.d(\col_addr_next[6]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[6]~q ),
	.prn(vcc));
defparam \col_addr_this[6] .is_wysiwyg = "true";
defparam \col_addr_this[6] .power_up = "low";

cycloneiii_lcell_comb \row_addr_next[7]~8 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[7]~8_combout ),
	.cout());
defparam \row_addr_next[7]~8 .lut_mask = 16'hEEEE;
defparam \row_addr_next[7]~8 .sum_lutc_input = "datac";

dffeas \row_addr_this[7] (
	.clk(clk),
	.d(\row_addr_next[7]~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[7]~q ),
	.prn(vcc));
defparam \row_addr_this[7] .is_wysiwyg = "true";
defparam \row_addr_this[7] .power_up = "low";

cycloneiii_lcell_comb \Selector29~0 (
	.dataa(\col_addr_this[6]~q ),
	.datab(\row_addr_this[7]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
defparam \Selector29~0 .lut_mask = 16'hACFF;
defparam \Selector29~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \col_addr_next[7]~7 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\col_addr_next[7]~7_combout ),
	.cout());
defparam \col_addr_next[7]~7 .lut_mask = 16'hEEEE;
defparam \col_addr_next[7]~7 .sum_lutc_input = "datac";

dffeas \col_addr_this[7] (
	.clk(clk),
	.d(\col_addr_next[7]~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\col_addr_this[7]~q ),
	.prn(vcc));
defparam \col_addr_this[7] .is_wysiwyg = "true";
defparam \col_addr_this[7] .power_up = "low";

dffeas \row_addr_this[8] (
	.clk(clk),
	.d(\row_addr_next[8]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[8]~q ),
	.prn(vcc));
defparam \row_addr_this[8] .is_wysiwyg = "true";
defparam \row_addr_this[8] .power_up = "low";

cycloneiii_lcell_comb \Selector28~0 (
	.dataa(\col_addr_this[7]~q ),
	.datab(\row_addr_this[8]~q ),
	.datac(\a[5]~600_combout ),
	.datad(\a[5]~614_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
defparam \Selector28~0 .lut_mask = 16'hACFF;
defparam \Selector28~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[9]~0 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[9]~0_combout ),
	.cout());
defparam \row_addr_next[9]~0 .lut_mask = 16'hEEEE;
defparam \row_addr_next[9]~0 .sum_lutc_input = "datac";

dffeas \row_addr_this[9] (
	.clk(clk),
	.d(\row_addr_next[9]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[9]~q ),
	.prn(vcc));
defparam \row_addr_this[9] .is_wysiwyg = "true";
defparam \row_addr_this[9] .power_up = "low";

cycloneiii_lcell_comb \Selector27~0 (
	.dataa(\a[0]~589_combout ),
	.datab(\row_addr_this[9]~q ),
	.datac(gnd),
	.datad(\a[0]~590_combout ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
defparam \Selector27~0 .lut_mask = 16'hEEFF;
defparam \Selector27~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \row_addr_next[10]~12 (
	.dataa(\in_buf|my_fifo|pipefull[0]~q ),
	.datab(\in_buf|my_fifo|pipe[0][20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\row_addr_next[10]~12_combout ),
	.cout());
defparam \row_addr_next[10]~12 .lut_mask = 16'hEEEE;
defparam \row_addr_next[10]~12 .sum_lutc_input = "datac";

dffeas \row_addr_this[10] (
	.clk(clk),
	.d(\row_addr_next[10]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[10]~q ),
	.prn(vcc));
defparam \row_addr_this[10] .is_wysiwyg = "true";
defparam \row_addr_this[10] .power_up = "low";

cycloneiii_lcell_comb \Selector26~1 (
	.dataa(\state.s_write~q ),
	.datab(\Selector5~6_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\p_main_fsm~154_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
defparam \Selector26~1 .lut_mask = 16'hFEFF;
defparam \Selector26~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector26~2 (
	.dataa(\Selector39~1_combout ),
	.datab(\Selector26~1_combout ),
	.datac(\Selector20~2_combout ),
	.datad(\p_main_fsm~170_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
defparam \Selector26~2 .lut_mask = 16'hFEFF;
defparam \Selector26~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~5 (
	.dataa(\state.s_holding~q ),
	.datab(\didnt_act~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
defparam \Selector5~5 .lut_mask = 16'hEEEE;
defparam \Selector5~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector26~0 (
	.dataa(\p_main_fsm~57_combout ),
	.datab(\Selector5~2_combout ),
	.datac(\Selector5~4_combout ),
	.datad(\Selector5~5_combout ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hBFFF;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector26~3 (
	.dataa(\Selector23~3_combout ),
	.datab(\row_addr_this[10]~q ),
	.datac(\Selector26~2_combout ),
	.datad(\Selector26~0_combout ),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
defparam \Selector26~3 .lut_mask = 16'hFEFF;
defparam \Selector26~3 .sum_lutc_input = "datac";

dffeas \row_addr_this[11] (
	.clk(clk),
	.d(\row_addr_next[11]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[11]~q ),
	.prn(vcc));
defparam \row_addr_this[11] .is_wysiwyg = "true";
defparam \row_addr_this[11] .power_up = "low";

cycloneiii_lcell_comb \Selector25~0 (
	.dataa(\a[0]~589_combout ),
	.datab(\row_addr_this[11]~q ),
	.datac(gnd),
	.datad(\a[0]~590_combout ),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
defparam \Selector25~0 .lut_mask = 16'hEEFF;
defparam \Selector25~0 .sum_lutc_input = "datac";

dffeas \row_addr_this[12] (
	.clk(clk),
	.d(\row_addr_next[12]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\accepted~q ),
	.q(\row_addr_this[12]~q ),
	.prn(vcc));
defparam \row_addr_this[12] .is_wysiwyg = "true";
defparam \row_addr_this[12] .power_up = "low";

cycloneiii_lcell_comb \Selector24~0 (
	.dataa(\a[0]~589_combout ),
	.datab(\row_addr_this[12]~q ),
	.datac(gnd),
	.datad(\a[0]~590_combout ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hEEFF;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~328 (
	.dataa(\bank_is_open~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\this_row_is_open~q ),
	.cin(gnd),
	.combout(\state~328_combout ),
	.cout());
defparam \state~328 .lut_mask = 16'hAAFF;
defparam \state~328 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~172 (
	.dataa(\am_writing~q ),
	.datab(\am_reading~q ),
	.datac(\finished_tras_all~q ),
	.datad(\Mux2~1_combout ),
	.cin(gnd),
	.combout(\p_main_fsm~172_combout ),
	.cout());
defparam \p_main_fsm~172 .lut_mask = 16'hEFFF;
defparam \p_main_fsm~172 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~141 (
	.dataa(\ba[1]~140_combout ),
	.datab(\state.s_idle~q ),
	.datac(\state~328_combout ),
	.datad(\p_main_fsm~172_combout ),
	.cin(gnd),
	.combout(\ba[1]~141_combout ),
	.cout());
defparam \ba[1]~141 .lut_mask = 16'hFEFF;
defparam \ba[1]~141 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~148 (
	.dataa(\ba[1]~147_combout ),
	.datab(\ba[1]~116_combout ),
	.datac(\read_req_this~q ),
	.datad(\state.s_write~q ),
	.cin(gnd),
	.combout(\ba[1]~148_combout ),
	.cout());
defparam \ba[1]~148 .lut_mask = 16'hFFFE;
defparam \ba[1]~148 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~149 (
	.dataa(\ba[1]~146_combout ),
	.datab(\ba[1]~148_combout ),
	.datac(\state.s_idle~q ),
	.datad(seq_ac_add_1t_ac_lat_internal),
	.cin(gnd),
	.combout(\ba[1]~149_combout ),
	.cout());
defparam \ba[1]~149 .lut_mask = 16'hFEFF;
defparam \ba[1]~149 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~150 (
	.dataa(\ba[1]~144_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ba[1]~149_combout ),
	.cin(gnd),
	.combout(\ba[1]~150_combout ),
	.cout());
defparam \ba[1]~150 .lut_mask = 16'hAAFF;
defparam \ba[1]~150 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~129 (
	.dataa(\size_last[1]~q ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\state.s_read~q ),
	.datad(\p_main_fsm~156_combout ),
	.cin(gnd),
	.combout(\ba[1]~129_combout ),
	.cout());
defparam \ba[1]~129 .lut_mask = 16'hFEFF;
defparam \ba[1]~129 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~151 (
	.dataa(\state.s_idle~q ),
	.datab(\bank_is_open~q ),
	.datac(\a[5]~575_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ba[1]~151_combout ),
	.cout());
defparam \ba[1]~151 .lut_mask = 16'hFEFE;
defparam \ba[1]~151 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~152 (
	.dataa(\ba[1]~123_combout ),
	.datab(\ba[1]~129_combout ),
	.datac(\ba[1]~151_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ba[1]~152_combout ),
	.cout());
defparam \ba[1]~152 .lut_mask = 16'hFEFE;
defparam \ba[1]~152 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~153 (
	.dataa(\ba[1]~135_combout ),
	.datab(\ba[1]~141_combout ),
	.datac(\ba[1]~150_combout ),
	.datad(\ba[1]~152_combout ),
	.cin(gnd),
	.combout(\ba[1]~153_combout ),
	.cout());
defparam \ba[1]~153 .lut_mask = 16'hEFFF;
defparam \ba[1]~153 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~156 (
	.dataa(\Selector5~3_combout ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\p_main_fsm~157_combout ),
	.datad(\wdata_burst_count[1]~51_combout ),
	.cin(gnd),
	.combout(\ba[1]~156_combout ),
	.cout());
defparam \ba[1]~156 .lut_mask = 16'hEFFF;
defparam \ba[1]~156 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~144 (
	.dataa(\ba[1]~142_combout ),
	.datab(\ba[1]~143_combout ),
	.datac(\bank_is_open~q ),
	.datad(\ba[1]~128_combout ),
	.cin(gnd),
	.combout(\ba[1]~144_combout ),
	.cout());
defparam \ba[1]~144 .lut_mask = 16'hEFFF;
defparam \ba[1]~144 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~157 (
	.dataa(\ba[1]~162_combout ),
	.datab(\ba[1]~156_combout ),
	.datac(\ba[1]~144_combout ),
	.datad(\ba[1]~149_combout ),
	.cin(gnd),
	.combout(\ba[1]~157_combout ),
	.cout());
defparam \ba[1]~157 .lut_mask = 16'hFFFE;
defparam \ba[1]~157 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~159 (
	.dataa(\state.s_read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state~333_combout ),
	.cin(gnd),
	.combout(\ba[1]~159_combout ),
	.cout());
defparam \ba[1]~159 .lut_mask = 16'hAAFF;
defparam \ba[1]~159 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~160 (
	.dataa(\state.s_write~q ),
	.datab(\state~328_combout ),
	.datac(\state.s_idle~q ),
	.datad(\p_main_fsm~19_combout ),
	.cin(gnd),
	.combout(\ba[1]~160_combout ),
	.cout());
defparam \ba[1]~160 .lut_mask = 16'hFEFF;
defparam \ba[1]~160 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ba[1]~161 (
	.dataa(\ba[1]~158_combout ),
	.datab(\ba[1]~159_combout ),
	.datac(\ba[1]~160_combout ),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\ba[1]~161_combout ),
	.cout());
defparam \ba[1]~161 .lut_mask = 16'hFEFF;
defparam \ba[1]~161 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector41~0 (
	.dataa(\bank_addr_this[0]~q ),
	.datab(\ba[1]~153_combout ),
	.datac(\ba[1]~157_combout ),
	.datad(\ba[1]~161_combout ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hEFFF;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector40~0 (
	.dataa(\bank_addr_this[1]~q ),
	.datab(\ba[1]~153_combout ),
	.datac(\ba[1]~157_combout ),
	.datad(\ba[1]~161_combout ),
	.cin(gnd),
	.combout(\Selector40~0_combout ),
	.cout());
defparam \Selector40~0 .lut_mask = 16'hEFFF;
defparam \Selector40~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~0 (
	.dataa(\p_main_fsm~19_combout ),
	.datab(\p_main_fsm~157_combout ),
	.datac(\p_main_fsm~154_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'h7FFF;
defparam \Selector18~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~1 (
	.dataa(\bank_is_open~q ),
	.datab(seq_ac_add_1t_ac_lat_internal),
	.datac(\p_main_fsm~154_combout ),
	.datad(\am_writing~q ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'hD8FF;
defparam \Selector18~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~3 (
	.dataa(\Selector18~2_combout ),
	.datab(\Mux2~1_combout ),
	.datac(\bank_is_open~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
defparam \Selector18~3 .lut_mask = 16'hFDFD;
defparam \Selector18~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~4 (
	.dataa(\state~331_combout ),
	.datab(\Selector18~0_combout ),
	.datac(\Selector18~1_combout ),
	.datad(\Selector18~3_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
defparam \Selector18~4 .lut_mask = 16'hEFFF;
defparam \Selector18~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \cs_n~63 (
	.dataa(\bank_is_open~q ),
	.datab(\Mux2~1_combout ),
	.datac(\p_main_fsm~171_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\cs_n~63_combout ),
	.cout());
defparam \cs_n~63 .lut_mask = 16'hBFFF;
defparam \cs_n~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~5 (
	.dataa(\p_main_fsm~156_combout ),
	.datab(\cs_n~63_combout ),
	.datac(\cs_n~64_combout ),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
defparam \Selector18~5 .lut_mask = 16'hFEFF;
defparam \Selector18~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector18~6 (
	.dataa(\Selector17~6_combout ),
	.datab(\Selector18~4_combout ),
	.datac(\Selector18~5_combout ),
	.datad(\Selector5~7_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
defparam \Selector18~6 .lut_mask = 16'hFF7F;
defparam \Selector18~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~7 (
	.dataa(\Selector19~9_combout ),
	.datab(\p_main_fsm~154_combout ),
	.datac(\Selector3~4_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector19~7_combout ),
	.cout());
defparam \Selector19~7 .lut_mask = 16'h8BFF;
defparam \Selector19~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~2 (
	.dataa(\am_writing~q ),
	.datab(\am_reading~q ),
	.datac(\am_reading_r~q ),
	.datad(\read_req_this~q ),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
defparam \Selector12~2 .lut_mask = 16'hFEFF;
defparam \Selector12~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector17~14 (
	.dataa(\new_req~49_combout ),
	.datab(\Selector12~2_combout ),
	.datac(gnd),
	.datad(\ba[1]~123_combout ),
	.cin(gnd),
	.combout(\Selector17~14_combout ),
	.cout());
defparam \Selector17~14 .lut_mask = 16'hEEFF;
defparam \Selector17~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~10 (
	.dataa(\rfsh_pending~q ),
	.datab(\refresh_in_progress~q ),
	.datac(\Selector17~14_combout ),
	.datad(\Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector19~10_combout ),
	.cout());
defparam \Selector19~10 .lut_mask = 16'hF7FF;
defparam \Selector19~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~168 (
	.dataa(\read_req_last~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\cs_addr_to_term[0]~q ),
	.cin(gnd),
	.combout(\p_main_fsm~168_combout ),
	.cout());
defparam \p_main_fsm~168 .lut_mask = 16'hAAFF;
defparam \p_main_fsm~168 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~0 (
	.dataa(\Selector43~1_combout ),
	.datab(\a[5]~574_combout ),
	.datac(\p_main_fsm~168_combout ),
	.datad(\p_main_fsm~158_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hEFFF;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~8 (
	.dataa(\Selector19~6_combout ),
	.datab(\Selector19~7_combout ),
	.datac(\Selector19~10_combout ),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(\Selector19~8_combout ),
	.cout());
defparam \Selector19~8 .lut_mask = 16'hFF7F;
defparam \Selector19~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~10 (
	.dataa(\Selector20~9_combout ),
	.datab(\state.s_holding~q ),
	.datac(\p_main_fsm~165_combout ),
	.datad(\Selector10~1_combout ),
	.cin(gnd),
	.combout(\Selector20~10_combout ),
	.cout());
defparam \Selector20~10 .lut_mask = 16'hFEFF;
defparam \Selector20~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~11 (
	.dataa(\Selector20~5_combout ),
	.datab(\state.s_write~q ),
	.datac(\p_main_fsm~105_combout ),
	.datad(\state~332_combout ),
	.cin(gnd),
	.combout(\Selector20~11_combout ),
	.cout());
defparam \Selector20~11 .lut_mask = 16'hFEFF;
defparam \Selector20~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector37~3 (
	.dataa(\state.s_read~q ),
	.datab(gnd),
	.datac(\size_last[1]~q ),
	.datad(\size_last[0]~q ),
	.cin(gnd),
	.combout(\Selector37~3_combout ),
	.cout());
defparam \Selector37~3 .lut_mask = 16'hAFFF;
defparam \Selector37~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~12 (
	.dataa(\Selector20~2_combout ),
	.datab(\state~328_combout ),
	.datac(\state.s_precharge~q ),
	.datad(\Selector37~3_combout ),
	.cin(gnd),
	.combout(\Selector20~12_combout ),
	.cout());
defparam \Selector20~12 .lut_mask = 16'hFFFB;
defparam \Selector20~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~13 (
	.dataa(\Selector20~3_combout ),
	.datab(\state.s_activate~q ),
	.datac(\Selector50~6_combout ),
	.datad(\Selector20~12_combout ),
	.cin(gnd),
	.combout(\Selector20~13_combout ),
	.cout());
defparam \Selector20~13 .lut_mask = 16'hFFEF;
defparam \Selector20~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~14 (
	.dataa(\Selector23~2_combout ),
	.datab(\bank_man|Equal8~0_combout ),
	.datac(\p_main_fsm~163_combout ),
	.datad(\Selector20~13_combout ),
	.cin(gnd),
	.combout(\Selector20~14_combout ),
	.cout());
defparam \Selector20~14 .lut_mask = 16'hFFFE;
defparam \Selector20~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~15 (
	.dataa(\Selector20~8_combout ),
	.datab(\Selector20~10_combout ),
	.datac(\Selector20~11_combout ),
	.datad(\Selector20~14_combout ),
	.cin(gnd),
	.combout(\Selector20~15_combout ),
	.cout());
defparam \Selector20~15 .lut_mask = 16'hFFFE;
defparam \Selector20~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~16 (
	.dataa(\state.s_reading~q ),
	.datab(\rdata_bcount_eq_1~q ),
	.datac(\didnt_term~q ),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\Selector20~16_combout ),
	.cout());
defparam \Selector20~16 .lut_mask = 16'hBFFF;
defparam \Selector20~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \p_main_fsm~173 (
	.dataa(\Mux2~1_combout ),
	.datab(\finished_tras~q ),
	.datac(\finished_tras_last~q ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\p_main_fsm~173_combout ),
	.cout());
defparam \p_main_fsm~173 .lut_mask = 16'h7FFF;
defparam \p_main_fsm~173 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~17 (
	.dataa(\Selector20~15_combout ),
	.datab(\Selector20~16_combout ),
	.datac(\Selector20~2_combout ),
	.datad(\p_main_fsm~173_combout ),
	.cin(gnd),
	.combout(\Selector20~17_combout ),
	.cout());
defparam \Selector20~17 .lut_mask = 16'h7FFF;
defparam \Selector20~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \control_wlat_r[0]~0 (
	.dataa(wd_lat_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_wlat_r[0]~0_combout ),
	.cout());
defparam \control_wlat_r[0]~0 .lut_mask = 16'h5555;
defparam \control_wlat_r[0]~0 .sum_lutc_input = "datac";

dffeas \control_wlat_r[1] (
	.clk(clk),
	.d(control_wlat[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\control_wlat_r[1]~q ),
	.prn(vcc));
defparam \control_wlat_r[1] .is_wysiwyg = "true";
defparam \control_wlat_r[1] .power_up = "low";

dffeas \control_wlat_r[4] (
	.clk(clk),
	.d(control_wlat[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\control_wlat_r[4]~q ),
	.prn(vcc));
defparam \control_wlat_r[4] .is_wysiwyg = "true";
defparam \control_wlat_r[4] .power_up = "low";

dffeas \control_wlat_r[3] (
	.clk(clk),
	.d(control_wlat[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\control_wlat_r[3]~q ),
	.prn(vcc));
defparam \control_wlat_r[3] .is_wysiwyg = "true";
defparam \control_wlat_r[3] .power_up = "low";

cycloneiii_lcell_comb \control_wlat_r[2]~1 (
	.dataa(wd_lat_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_wlat_r[2]~1_combout ),
	.cout());
defparam \control_wlat_r[2]~1 .lut_mask = 16'h5555;
defparam \control_wlat_r[2]~1 .sum_lutc_input = "datac";

dffeas \control_wlat_r[2] (
	.clk(clk),
	.d(\control_wlat_r[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\control_wlat_r[2]~q ),
	.prn(vcc));
defparam \control_wlat_r[2] .is_wysiwyg = "true";
defparam \control_wlat_r[2] .power_up = "low";

dffeas fifo_rdreq_cas4(
	.clk(clk),
	.d(\doing_wr_cl_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_rdreq_cas4~q ),
	.prn(vcc));
defparam fifo_rdreq_cas4.is_wysiwyg = "true";
defparam fifo_rdreq_cas4.power_up = "low";

dffeas fifo_rdreq_cas5(
	.clk(clk),
	.d(\fifo_rdreq_cas4~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_rdreq_cas5~q ),
	.prn(vcc));
defparam fifo_rdreq_cas5.is_wysiwyg = "true";
defparam fifo_rdreq_cas5.power_up = "low";

cycloneiii_lcell_comb \control_doing_wr~2 (
	.dataa(control_wlat_r_0),
	.datab(control_doing_wr),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_doing_wr~2_combout ),
	.cout());
defparam \control_doing_wr~2 .lut_mask = 16'hEEEE;
defparam \control_doing_wr~2 .sum_lutc_input = "datac";

dffeas fifo_rdreq_cas6(
	.clk(clk),
	.d(\fifo_rdreq_cas5~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_rdreq_cas6~q ),
	.prn(vcc));
defparam fifo_rdreq_cas6.is_wysiwyg = "true";
defparam fifo_rdreq_cas6.power_up = "low";

cycloneiii_lcell_comb \LessThan6~0 (
	.dataa(\dqs_must_keep_toggling[2]~q ),
	.datab(\dqs_must_keep_toggling[1]~q ),
	.datac(\dqs_must_keep_toggling[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan6~0_combout ),
	.cout());
defparam \LessThan6~0 .lut_mask = 16'hFEFE;
defparam \LessThan6~0 .sum_lutc_input = "datac";

dffeas dqs_brst_odd_dtt(
	.clk(clk),
	.d(\LessThan6~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_brst_odd_dtt~q ),
	.prn(vcc));
defparam dqs_brst_odd_dtt.is_wysiwyg = "true";
defparam dqs_brst_odd_dtt.power_up = "low";

endmodule

module altera_ddr_auk_ddr_hp_avalon_if (
	pipefull_3,
	clk,
	local_be,
	local_wdata,
	seq_ac_add_1t_ac_lat_internal,
	reset_phy_clk_1x_n,
	control_doing_wr,
	control_doing_wr1,
	local_write_req,
	avalon_be,
	avalon_wdata)/* synthesis synthesis_greybox=1 */;
input 	pipefull_3;
input 	clk;
output 	[3:0] local_be;
output 	[31:0] local_wdata;
input 	seq_ac_add_1t_ac_lat_internal;
input 	reset_phy_clk_1x_n;
input 	control_doing_wr;
input 	control_doing_wr1;
input 	local_write_req;
input 	[3:0] avalon_be;
input 	[31:0] avalon_wdata;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_scfifo_1 wfifo(
	.pipefull_3(pipefull_3),
	.clock(clk),
	.q({local_be[3],local_be[2],local_be[1],local_be[0],local_wdata[31],local_wdata[30],local_wdata[29],local_wdata[28],local_wdata[27],local_wdata[26],local_wdata[25],local_wdata[24],local_wdata[23],local_wdata[22],local_wdata[21],local_wdata[20],local_wdata[19],local_wdata[18],local_wdata[17],local_wdata[16],local_wdata[15],local_wdata[14],local_wdata[13],local_wdata[12],
local_wdata[11],local_wdata[10],local_wdata[9],local_wdata[8],local_wdata[7],local_wdata[6],local_wdata[5],local_wdata[4],local_wdata[3],local_wdata[2],local_wdata[1],local_wdata[0]}),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_wr(control_doing_wr),
	.control_doing_wr1(control_doing_wr1),
	.local_write_req(local_write_req),
	.data({avalon_be[3],avalon_be[2],avalon_be[1],avalon_be[0],avalon_wdata[31],avalon_wdata[30],avalon_wdata[29],avalon_wdata[28],avalon_wdata[27],avalon_wdata[26],avalon_wdata[25],avalon_wdata[24],avalon_wdata[23],avalon_wdata[22],avalon_wdata[21],avalon_wdata[20],avalon_wdata[19],avalon_wdata[18],avalon_wdata[17],avalon_wdata[16],avalon_wdata[15],avalon_wdata[14],
avalon_wdata[13],avalon_wdata[12],avalon_wdata[11],avalon_wdata[10],avalon_wdata[9],avalon_wdata[8],avalon_wdata[7],avalon_wdata[6],avalon_wdata[5],avalon_wdata[4],avalon_wdata[3],avalon_wdata[2],avalon_wdata[1],avalon_wdata[0]}));

endmodule

module altera_ddr_scfifo_1 (
	pipefull_3,
	clock,
	q,
	seq_ac_add_1t_ac_lat_internal,
	reset_phy_clk_1x_n,
	control_doing_wr,
	control_doing_wr1,
	local_write_req,
	data)/* synthesis synthesis_greybox=1 */;
input 	pipefull_3;
input 	clock;
output 	[35:0] q;
input 	seq_ac_add_1t_ac_lat_internal;
input 	reset_phy_clk_1x_n;
input 	control_doing_wr;
input 	control_doing_wr1;
input 	local_write_req;
input 	[35:0] data;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_scfifo_jve1 auto_generated(
	.pipefull_3(pipefull_3),
	.clock(clock),
	.q({q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_wr(control_doing_wr),
	.control_doing_wr1(control_doing_wr1),
	.local_write_req(local_write_req),
	.data({data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module altera_ddr_scfifo_jve1 (
	pipefull_3,
	clock,
	q,
	seq_ac_add_1t_ac_lat_internal,
	reset_phy_clk_1x_n,
	control_doing_wr,
	control_doing_wr1,
	local_write_req,
	data)/* synthesis synthesis_greybox=1 */;
input 	pipefull_3;
input 	clock;
output 	[35:0] q;
input 	seq_ac_add_1t_ac_lat_internal;
input 	reset_phy_clk_1x_n;
input 	control_doing_wr;
input 	control_doing_wr1;
input 	local_write_req;
input 	[35:0] data;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_a_dpfifo_kg71 dpfifo(
	.pipefull_3(pipefull_3),
	.clock(clock),
	.q({q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_wr(control_doing_wr),
	.control_doing_wr1(control_doing_wr1),
	.local_write_req(local_write_req),
	.data({data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module altera_ddr_a_dpfifo_kg71 (
	pipefull_3,
	clock,
	q,
	seq_ac_add_1t_ac_lat_internal,
	reset_phy_clk_1x_n,
	control_doing_wr,
	control_doing_wr1,
	local_write_req,
	data)/* synthesis synthesis_greybox=1 */;
input 	pipefull_3;
input 	clock;
output 	[35:0] q;
input 	seq_ac_add_1t_ac_lat_internal;
input 	reset_phy_clk_1x_n;
input 	control_doing_wr;
input 	control_doing_wr1;
input 	local_write_req;
input 	[35:0] data;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \full_dff~q ;
wire \valid_wreq~combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \low_addressa[0]~q ;
wire \empty_dff~q ;
wire \valid_rreq~combout ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~10_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~11_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~12_combout ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~13_combout ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~14_combout ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \_~63_combout ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \_~64_combout ;
wire \_~65_combout ;
wire \usedw_is_1_dff~q ;
wire \usedw_is_0_dff~q ;
wire \_~41_combout ;
wire \usedw_is_2_dff~q ;
wire \usedw_will_be_1~2_combout ;
wire \_~45_combout ;
wire \_~0_combout ;
wire \_~31_combout ;
wire \_~7_combout ;
wire \usedw_will_be_1~1_combout ;
wire \_~66_combout ;
wire \usedw_will_be_2~2_combout ;
wire \usedw_will_be_2~1_combout ;
wire \rd_ptr_lsb~3_combout ;


altera_ddr_altsyncram_1ea1 FIFOram(
	.clock0(clock),
	.q_b({q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren_a(\valid_wreq~combout ),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[4]~14_combout ,\ram_read_address[3]~13_combout ,\ram_read_address[2]~12_combout ,\ram_read_address[1]~11_combout ,\ram_read_address[0]~10_combout }),
	.data_a({data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

altera_ddr_cntr_mmb rd_ptr_msb(
	.clock(clock),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	._(\_~31_combout ));

altera_ddr_cntr_3n7 usedw_counter(
	.clock(clock),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.updown(\valid_wreq~combout ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	._(\_~7_combout ));

altera_ddr_cntr_nmb wr_ptr(
	.clock(clock),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.valid_wreq(\valid_wreq~combout ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ));

dffeas full_dff(
	.clk(clock),
	.d(\_~65_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneiii_lcell_comb valid_wreq(
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(local_write_req),
	.datac(pipefull_3),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~combout ),
	.cout());
defparam valid_wreq.lut_mask = 16'hEFFF;
defparam valid_wreq.sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~10_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas empty_dff(
	.clk(clock),
	.d(\_~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneiii_lcell_comb valid_rreq(
	.dataa(\empty_dff~q ),
	.datab(control_doing_wr),
	.datac(control_doing_wr1),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_rreq~combout ),
	.cout());
defparam valid_rreq.lut_mask = 16'hFEFE;
defparam valid_rreq.sum_lutc_input = "datac";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~3_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_rreq~combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneiii_lcell_comb \ram_read_address[0]~10 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~10_combout ),
	.cout());
defparam \ram_read_address[0]~10 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~10 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[1]~11 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~11_combout ),
	.cout());
defparam \ram_read_address[1]~11 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~11 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[2]~12 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~12_combout ),
	.cout());
defparam \ram_read_address[2]~12 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~12 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\ram_read_address[3]~13_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[3]~13 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~13_combout ),
	.cout());
defparam \ram_read_address[3]~13 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~13 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\ram_read_address[4]~14_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneiii_lcell_comb \ram_read_address[4]~14 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~14_combout ),
	.cout());
defparam \ram_read_address[4]~14 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~63 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~63_combout ),
	.cout());
defparam \_~63 .lut_mask = 16'hEEEE;
defparam \_~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~64 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~63_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~64_combout ),
	.cout());
defparam \_~64 .lut_mask = 16'hFFFE;
defparam \_~64 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~65 (
	.dataa(\full_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(\_~64_combout ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\_~65_combout ),
	.cout());
defparam \_~65 .lut_mask = 16'hFEFF;
defparam \_~65 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\_~41_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneiii_lcell_comb \_~41 (
	.dataa(\valid_rreq~combout ),
	.datab(\usedw_is_1_dff~q ),
	.datac(\valid_wreq~combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\_~41_combout ),
	.cout());
defparam \_~41 .lut_mask = 16'hFF7B;
defparam \_~41 .sum_lutc_input = "datac";

dffeas usedw_is_2_dff(
	.clk(clock),
	.d(\usedw_will_be_2~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_2_dff~q ),
	.prn(vcc));
defparam usedw_is_2_dff.is_wysiwyg = "true";
defparam usedw_is_2_dff.power_up = "low";

cycloneiii_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(\valid_rreq~combout ),
	.datac(\usedw_is_0_dff~q ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFEF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~45 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(\valid_rreq~combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\_~45_combout ),
	.cout());
defparam \_~45 .lut_mask = 16'hBEBE;
defparam \_~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~0 (
	.dataa(\_~41_combout ),
	.datab(\valid_wreq~combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(\_~45_combout ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hBFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~31 (
	.dataa(\empty_dff~q ),
	.datab(control_doing_wr),
	.datac(control_doing_wr1),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\_~31_combout ),
	.cout());
defparam \_~31 .lut_mask = 16'hFEFF;
defparam \_~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~7 (
	.dataa(control_doing_wr),
	.datab(control_doing_wr1),
	.datac(\valid_wreq~combout ),
	.datad(\empty_dff~q ),
	.cin(gnd),
	.combout(\_~7_combout ),
	.cout());
defparam \_~7 .lut_mask = 16'h6996;
defparam \_~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_will_be_1~2_combout ),
	.datab(\usedw_is_1_dff~q ),
	.datac(\valid_wreq~combout ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hEFFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \_~66 (
	.dataa(\_~63_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~66_combout ),
	.cout());
defparam \_~66 .lut_mask = 16'hBFFF;
defparam \_~66 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \usedw_will_be_2~2 (
	.dataa(\usedw_is_2_dff~q ),
	.datab(\valid_rreq~combout ),
	.datac(\_~66_combout ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_2~2_combout ),
	.cout());
defparam \usedw_will_be_2~2 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_2~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \usedw_will_be_2~1 (
	.dataa(\usedw_will_be_2~2_combout ),
	.datab(\valid_wreq~combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_2~1_combout ),
	.cout());
defparam \usedw_will_be_2~1 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ptr_lsb~3 (
	.dataa(\rd_ptr_lsb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ptr_lsb~3_combout ),
	.cout());
defparam \rd_ptr_lsb~3 .lut_mask = 16'h5555;
defparam \rd_ptr_lsb~3 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altsyncram_1ea1 (
	clock0,
	q_b,
	wren_a,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[35:0] q_b;
input 	wren_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	[35:0] data_a;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;


wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a34(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus));
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 5;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 31;
defparam ram_block1a34.port_a_logical_ram_depth = 32;
defparam ram_block1a34.port_a_logical_ram_width = 36;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock0";
defparam ram_block1a34.port_b_address_width = 5;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "none";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 31;
defparam ram_block1a34.port_b_logical_ram_depth = 32;
defparam ram_block1a34.port_b_logical_ram_width = 36;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock0";
defparam ram_block1a34.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a32(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus));
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 5;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 31;
defparam ram_block1a32.port_a_logical_ram_depth = 32;
defparam ram_block1a32.port_a_logical_ram_width = 36;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock0";
defparam ram_block1a32.port_b_address_width = 5;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "none";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 31;
defparam ram_block1a32.port_b_logical_ram_depth = 32;
defparam ram_block1a32.port_b_logical_ram_width = 36;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock0";
defparam ram_block1a32.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a35(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus));
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 5;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 31;
defparam ram_block1a35.port_a_logical_ram_depth = 32;
defparam ram_block1a35.port_a_logical_ram_width = 36;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock0";
defparam ram_block1a35.port_b_address_width = 5;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "none";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 31;
defparam ram_block1a35.port_b_logical_ram_depth = 32;
defparam ram_block1a35.port_b_logical_ram_width = 36;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock0";
defparam ram_block1a35.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a33(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus));
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 5;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 31;
defparam ram_block1a33.port_a_logical_ram_depth = 32;
defparam ram_block1a33.port_a_logical_ram_width = 36;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock0";
defparam ram_block1a33.port_b_address_width = 5;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "none";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 31;
defparam ram_block1a33.port_b_logical_ram_depth = 32;
defparam ram_block1a33.port_b_logical_ram_width = 36;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock0";
defparam ram_block1a33.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 36;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 36;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 36;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 36;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 36;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 36;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 36;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 36;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 36;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 36;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 36;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 36;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 36;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 36;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 36;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 36;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 36;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 36;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 36;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 36;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 36;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 36;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 36;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 36;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 36;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 36;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 36;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 36;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 36;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 36;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 36;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 36;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 36;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 36;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 36;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 36;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 36;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 36;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 36;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 36;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 36;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 36;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 36;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 36;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 36;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 36;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 36;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 36;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 36;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 36;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 36;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 36;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 36;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 36;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 36;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 36;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 36;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 36;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 36;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 36;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 36;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 36;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_auk_ddr_hp_controller_wrapper:altera_ddr_auk_ddr_hp_controller_wrapper_inst|auk_ddr_hp_controller:auk_ddr_hp_controller_inst|auk_ddr_hp_avalon_if:\\g_local_avalon_if:av_if|scfifo:wfifo|scfifo_jve1:auto_generated|a_dpfifo_kg71:dpfifo|altsyncram_1ea1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 36;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 36;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

endmodule

module altera_ddr_cntr_3n7 (
	clock,
	reset_phy_clk_1x_n,
	updown,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	_)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	reset_phy_clk_1x_n;
input 	updown;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	_;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module altera_ddr_cntr_mmb (
	clock,
	reset_phy_clk_1x_n,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	_)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	reset_phy_clk_1x_n;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	_;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module altera_ddr_cntr_nmb (
	clock,
	reset_phy_clk_1x_n,
	valid_wreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	reset_phy_clk_1x_n;
input 	valid_wreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_wreq),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_wreq),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_wreq),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_wreq),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(valid_wreq),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneiii_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneiii_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module altera_ddr_auk_ddr_hp_bank_details (
	clk,
	reset_n,
	Equal8,
	doing_act,
	in_this_bank,
	doing_pch_all,
	doing_pch,
	row_mux_sel_next_1,
	row_mux_sel_next_0,
	Mux11,
	Mux3,
	Mux8,
	Mux2,
	Mux9,
	Mux4,
	Mux12,
	Mux7,
	Mux5,
	Mux6,
	Mux10,
	Mux1,
	Mux0,
	Mux13,
	row_addr_this_0,
	row_addr_this_1,
	row_addr_this_2,
	row_addr_this_3,
	row_addr_this_4,
	row_addr_this_5,
	row_addr_this_6,
	row_addr_this_7,
	row_addr_this_8,
	row_addr_this_9,
	row_addr_this_10,
	row_addr_this_11,
	row_addr_this_12)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
output 	Equal8;
input 	doing_act;
input 	[2:0] in_this_bank;
input 	doing_pch_all;
input 	doing_pch;
input 	row_mux_sel_next_1;
input 	row_mux_sel_next_0;
output 	Mux11;
output 	Mux3;
output 	Mux8;
output 	Mux2;
output 	Mux9;
output 	Mux4;
output 	Mux12;
output 	Mux7;
output 	Mux5;
output 	Mux6;
output 	Mux10;
output 	Mux1;
output 	Mux0;
output 	Mux13;
input 	row_addr_this_0;
input 	row_addr_this_1;
input 	row_addr_this_2;
input 	row_addr_this_3;
input 	row_addr_this_4;
input 	row_addr_this_5;
input 	row_addr_this_6;
input 	row_addr_this_7;
input 	row_addr_this_8;
input 	row_addr_this_9;
input 	row_addr_this_10;
input 	row_addr_this_11;
input 	row_addr_this_12;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \in_this_bank_r[0]~q ;
wire \in_this_bank_r[1]~q ;
wire \bank_is_open[3]~32_combout ;
wire \bank_is_open[3]~33_combout ;
wire \bank_is_open[3]~q ;
wire \bank_is_open[2]~34_combout ;
wire \bank_is_open[2]~35_combout ;
wire \bank_is_open[2]~q ;
wire \bank_is_open[1]~36_combout ;
wire \bank_is_open[1]~37_combout ;
wire \bank_is_open[1]~q ;
wire \bank_is_open[0]~38_combout ;
wire \bank_is_open[0]~39_combout ;
wire \bank_is_open[0]~q ;
wire \openrows~416_combout ;
wire \openrows[1][8]~417_combout ;
wire \openrows[2][11]~418_combout ;
wire \openrows[2][1]~q ;
wire \openrows[1][8]~419_combout ;
wire \openrows[1][1]~q ;
wire \openrows[0][2]~420_combout ;
wire \openrows[0][1]~q ;
wire \Mux11~0_combout ;
wire \openrows[3][5]~421_combout ;
wire \openrows[3][1]~q ;
wire \openrows~422_combout ;
wire \openrows[2][9]~q ;
wire \openrows[1][9]~q ;
wire \openrows[0][9]~q ;
wire \Mux3~0_combout ;
wire \openrows[3][9]~q ;
wire \openrows~423_combout ;
wire \openrows[1][4]~q ;
wire \openrows[2][4]~q ;
wire \openrows[0][4]~q ;
wire \Mux8~0_combout ;
wire \openrows[3][4]~q ;
wire \openrows~424_combout ;
wire \openrows[1][10]~q ;
wire \openrows[2][10]~q ;
wire \openrows[0][10]~q ;
wire \Mux2~0_combout ;
wire \openrows[3][10]~q ;
wire \openrows~425_combout ;
wire \openrows[2][3]~q ;
wire \openrows[1][3]~q ;
wire \openrows[0][3]~q ;
wire \Mux9~0_combout ;
wire \openrows[3][3]~q ;
wire \openrows~426_combout ;
wire \openrows[1][8]~q ;
wire \openrows[2][8]~q ;
wire \openrows[0][8]~q ;
wire \Mux4~0_combout ;
wire \openrows[3][8]~q ;
wire \openrows~427_combout ;
wire \openrows[1][0]~q ;
wire \openrows[2][0]~q ;
wire \openrows[0][0]~q ;
wire \Mux12~0_combout ;
wire \openrows[3][0]~q ;
wire \openrows~428_combout ;
wire \openrows[2][5]~q ;
wire \openrows[1][5]~q ;
wire \openrows[0][5]~q ;
wire \Mux7~0_combout ;
wire \openrows[3][5]~q ;
wire \openrows~429_combout ;
wire \openrows[2][7]~q ;
wire \openrows[1][7]~q ;
wire \openrows[0][7]~q ;
wire \Mux5~0_combout ;
wire \openrows[3][7]~q ;
wire \openrows~430_combout ;
wire \openrows[1][6]~q ;
wire \openrows[2][6]~q ;
wire \openrows[0][6]~q ;
wire \Mux6~0_combout ;
wire \openrows[3][6]~q ;
wire \openrows~431_combout ;
wire \openrows[1][2]~q ;
wire \openrows[2][2]~q ;
wire \openrows[0][2]~q ;
wire \Mux10~0_combout ;
wire \openrows[3][2]~q ;
wire \openrows~432_combout ;
wire \openrows[2][11]~q ;
wire \openrows[1][11]~q ;
wire \openrows[0][11]~q ;
wire \Mux1~0_combout ;
wire \openrows[3][11]~q ;
wire \openrows~433_combout ;
wire \openrows[1][12]~q ;
wire \openrows[2][12]~q ;
wire \openrows[0][12]~q ;
wire \Mux0~0_combout ;
wire \openrows[3][12]~q ;
wire \Mux13~0_combout ;


cycloneiii_lcell_comb \Equal8~0 (
	.dataa(\bank_is_open[3]~q ),
	.datab(\bank_is_open[2]~q ),
	.datac(\bank_is_open[1]~q ),
	.datad(\bank_is_open[0]~q ),
	.cin(gnd),
	.combout(Equal8),
	.cout());
defparam \Equal8~0 .lut_mask = 16'h7FFF;
defparam \Equal8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux11~1 (
	.dataa(\openrows[2][1]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux11~0_combout ),
	.datad(\openrows[3][1]~q ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
defparam \Mux11~1 .lut_mask = 16'hFFBE;
defparam \Mux11~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux3~1 (
	.dataa(\openrows[2][9]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux3~0_combout ),
	.datad(\openrows[3][9]~q ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux8~1 (
	.dataa(\openrows[1][4]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux8~0_combout ),
	.datad(\openrows[3][4]~q ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hFFBE;
defparam \Mux8~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux2~1 (
	.dataa(\openrows[1][10]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux2~0_combout ),
	.datad(\openrows[3][10]~q ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux9~1 (
	.dataa(\openrows[2][3]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux9~0_combout ),
	.datad(\openrows[3][3]~q ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hFFBE;
defparam \Mux9~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux4~1 (
	.dataa(\openrows[1][8]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux4~0_combout ),
	.datad(\openrows[3][8]~q ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFFBE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux12~1 (
	.dataa(\openrows[1][0]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux12~0_combout ),
	.datad(\openrows[3][0]~q ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
defparam \Mux12~1 .lut_mask = 16'hFFBE;
defparam \Mux12~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux7~1 (
	.dataa(\openrows[2][5]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux7~0_combout ),
	.datad(\openrows[3][5]~q ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hFFBE;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux5~1 (
	.dataa(\openrows[2][7]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux5~0_combout ),
	.datad(\openrows[3][7]~q ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFFBE;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux6~1 (
	.dataa(\openrows[1][6]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux6~0_combout ),
	.datad(\openrows[3][6]~q ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hFFBE;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux10~1 (
	.dataa(\openrows[1][2]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux10~0_combout ),
	.datad(\openrows[3][2]~q ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
defparam \Mux10~1 .lut_mask = 16'hFFBE;
defparam \Mux10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(\openrows[2][11]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux1~0_combout ),
	.datad(\openrows[3][11]~q ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(\openrows[1][12]~q ),
	.datab(row_mux_sel_next_0),
	.datac(\Mux0~0_combout ),
	.datad(\openrows[3][12]~q ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux13~1 (
	.dataa(\bank_is_open[2]~q ),
	.datab(row_mux_sel_next_1),
	.datac(\Mux13~0_combout ),
	.datad(\bank_is_open[3]~q ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
defparam \Mux13~1 .lut_mask = 16'hFFBE;
defparam \Mux13~1 .sum_lutc_input = "datac";

dffeas \in_this_bank_r[0] (
	.clk(clk),
	.d(in_this_bank[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset_n),
	.q(\in_this_bank_r[0]~q ),
	.prn(vcc));
defparam \in_this_bank_r[0] .is_wysiwyg = "true";
defparam \in_this_bank_r[0] .power_up = "low";

dffeas \in_this_bank_r[1] (
	.clk(clk),
	.d(in_this_bank[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset_n),
	.q(\in_this_bank_r[1]~q ),
	.prn(vcc));
defparam \in_this_bank_r[1] .is_wysiwyg = "true";
defparam \in_this_bank_r[1] .power_up = "low";

cycloneiii_lcell_comb \bank_is_open[3]~32 (
	.dataa(doing_pch),
	.datab(\in_this_bank_r[0]~q ),
	.datac(\in_this_bank_r[1]~q ),
	.datad(doing_act),
	.cin(gnd),
	.combout(\bank_is_open[3]~32_combout ),
	.cout());
defparam \bank_is_open[3]~32 .lut_mask = 16'hFFFE;
defparam \bank_is_open[3]~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \bank_is_open[3]~33 (
	.dataa(\bank_is_open[3]~q ),
	.datab(doing_pch_all),
	.datac(doing_pch),
	.datad(\bank_is_open[3]~32_combout ),
	.cin(gnd),
	.combout(\bank_is_open[3]~33_combout ),
	.cout());
defparam \bank_is_open[3]~33 .lut_mask = 16'hAF3F;
defparam \bank_is_open[3]~33 .sum_lutc_input = "datac";

dffeas \bank_is_open[3] (
	.clk(clk),
	.d(\bank_is_open[3]~33_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bank_is_open[3]~q ),
	.prn(vcc));
defparam \bank_is_open[3] .is_wysiwyg = "true";
defparam \bank_is_open[3] .power_up = "low";

cycloneiii_lcell_comb \bank_is_open[2]~34 (
	.dataa(doing_pch),
	.datab(\in_this_bank_r[0]~q ),
	.datac(\in_this_bank_r[1]~q ),
	.datad(doing_act),
	.cin(gnd),
	.combout(\bank_is_open[2]~34_combout ),
	.cout());
defparam \bank_is_open[2]~34 .lut_mask = 16'hFFFB;
defparam \bank_is_open[2]~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \bank_is_open[2]~35 (
	.dataa(\bank_is_open[2]~q ),
	.datab(doing_pch_all),
	.datac(doing_pch),
	.datad(\bank_is_open[2]~34_combout ),
	.cin(gnd),
	.combout(\bank_is_open[2]~35_combout ),
	.cout());
defparam \bank_is_open[2]~35 .lut_mask = 16'hAF3F;
defparam \bank_is_open[2]~35 .sum_lutc_input = "datac";

dffeas \bank_is_open[2] (
	.clk(clk),
	.d(\bank_is_open[2]~35_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bank_is_open[2]~q ),
	.prn(vcc));
defparam \bank_is_open[2] .is_wysiwyg = "true";
defparam \bank_is_open[2] .power_up = "low";

cycloneiii_lcell_comb \bank_is_open[1]~36 (
	.dataa(doing_pch),
	.datab(\in_this_bank_r[1]~q ),
	.datac(\in_this_bank_r[0]~q ),
	.datad(doing_act),
	.cin(gnd),
	.combout(\bank_is_open[1]~36_combout ),
	.cout());
defparam \bank_is_open[1]~36 .lut_mask = 16'hFFFB;
defparam \bank_is_open[1]~36 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \bank_is_open[1]~37 (
	.dataa(\bank_is_open[1]~q ),
	.datab(doing_pch_all),
	.datac(doing_pch),
	.datad(\bank_is_open[1]~36_combout ),
	.cin(gnd),
	.combout(\bank_is_open[1]~37_combout ),
	.cout());
defparam \bank_is_open[1]~37 .lut_mask = 16'hAF3F;
defparam \bank_is_open[1]~37 .sum_lutc_input = "datac";

dffeas \bank_is_open[1] (
	.clk(clk),
	.d(\bank_is_open[1]~37_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bank_is_open[1]~q ),
	.prn(vcc));
defparam \bank_is_open[1] .is_wysiwyg = "true";
defparam \bank_is_open[1] .power_up = "low";

cycloneiii_lcell_comb \bank_is_open[0]~38 (
	.dataa(doing_pch),
	.datab(\in_this_bank_r[0]~q ),
	.datac(\in_this_bank_r[1]~q ),
	.datad(doing_act),
	.cin(gnd),
	.combout(\bank_is_open[0]~38_combout ),
	.cout());
defparam \bank_is_open[0]~38 .lut_mask = 16'hFFBF;
defparam \bank_is_open[0]~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \bank_is_open[0]~39 (
	.dataa(\bank_is_open[0]~q ),
	.datab(doing_pch_all),
	.datac(doing_pch),
	.datad(\bank_is_open[0]~38_combout ),
	.cin(gnd),
	.combout(\bank_is_open[0]~39_combout ),
	.cout());
defparam \bank_is_open[0]~39 .lut_mask = 16'hAF3F;
defparam \bank_is_open[0]~39 .sum_lutc_input = "datac";

dffeas \bank_is_open[0] (
	.clk(clk),
	.d(\bank_is_open[0]~39_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bank_is_open[0]~q ),
	.prn(vcc));
defparam \bank_is_open[0] .is_wysiwyg = "true";
defparam \bank_is_open[0] .power_up = "low";

cycloneiii_lcell_comb \openrows~416 (
	.dataa(row_addr_this_1),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~416_combout ),
	.cout());
defparam \openrows~416 .lut_mask = 16'hAFFF;
defparam \openrows~416 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \openrows[1][8]~417 (
	.dataa(gnd),
	.datab(gnd),
	.datac(doing_act),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows[1][8]~417_combout ),
	.cout());
defparam \openrows[1][8]~417 .lut_mask = 16'h0FFF;
defparam \openrows[1][8]~417 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \openrows[2][11]~418 (
	.dataa(\in_this_bank_r[0]~q ),
	.datab(\openrows[1][8]~417_combout ),
	.datac(\in_this_bank_r[1]~q ),
	.datad(doing_pch_all),
	.cin(gnd),
	.combout(\openrows[2][11]~418_combout ),
	.cout());
defparam \openrows[2][11]~418 .lut_mask = 16'hFFF7;
defparam \openrows[2][11]~418 .sum_lutc_input = "datac";

dffeas \openrows[2][1] (
	.clk(clk),
	.d(\openrows~416_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][1]~q ),
	.prn(vcc));
defparam \openrows[2][1] .is_wysiwyg = "true";
defparam \openrows[2][1] .power_up = "low";

cycloneiii_lcell_comb \openrows[1][8]~419 (
	.dataa(\in_this_bank_r[1]~q ),
	.datab(\openrows[1][8]~417_combout ),
	.datac(\in_this_bank_r[0]~q ),
	.datad(doing_pch_all),
	.cin(gnd),
	.combout(\openrows[1][8]~419_combout ),
	.cout());
defparam \openrows[1][8]~419 .lut_mask = 16'hFFF7;
defparam \openrows[1][8]~419 .sum_lutc_input = "datac";

dffeas \openrows[1][1] (
	.clk(clk),
	.d(\openrows~416_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][1]~q ),
	.prn(vcc));
defparam \openrows[1][1] .is_wysiwyg = "true";
defparam \openrows[1][1] .power_up = "low";

cycloneiii_lcell_comb \openrows[0][2]~420 (
	.dataa(\in_this_bank_r[0]~q ),
	.datab(\in_this_bank_r[1]~q ),
	.datac(\openrows[1][8]~417_combout ),
	.datad(doing_pch_all),
	.cin(gnd),
	.combout(\openrows[0][2]~420_combout ),
	.cout());
defparam \openrows[0][2]~420 .lut_mask = 16'hFF7F;
defparam \openrows[0][2]~420 .sum_lutc_input = "datac";

dffeas \openrows[0][1] (
	.clk(clk),
	.d(\openrows~416_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][1]~q ),
	.prn(vcc));
defparam \openrows[0][1] .is_wysiwyg = "true";
defparam \openrows[0][1] .power_up = "low";

cycloneiii_lcell_comb \Mux11~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][1]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][1]~q ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hFFDE;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \openrows[3][5]~421 (
	.dataa(\openrows[1][8]~417_combout ),
	.datab(\in_this_bank_r[0]~q ),
	.datac(\in_this_bank_r[1]~q ),
	.datad(doing_pch_all),
	.cin(gnd),
	.combout(\openrows[3][5]~421_combout ),
	.cout());
defparam \openrows[3][5]~421 .lut_mask = 16'hFFFD;
defparam \openrows[3][5]~421 .sum_lutc_input = "datac";

dffeas \openrows[3][1] (
	.clk(clk),
	.d(\openrows~416_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][1]~q ),
	.prn(vcc));
defparam \openrows[3][1] .is_wysiwyg = "true";
defparam \openrows[3][1] .power_up = "low";

cycloneiii_lcell_comb \openrows~422 (
	.dataa(row_addr_this_9),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~422_combout ),
	.cout());
defparam \openrows~422 .lut_mask = 16'hAFFF;
defparam \openrows~422 .sum_lutc_input = "datac";

dffeas \openrows[2][9] (
	.clk(clk),
	.d(\openrows~422_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][9]~q ),
	.prn(vcc));
defparam \openrows[2][9] .is_wysiwyg = "true";
defparam \openrows[2][9] .power_up = "low";

dffeas \openrows[1][9] (
	.clk(clk),
	.d(\openrows~422_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][9]~q ),
	.prn(vcc));
defparam \openrows[1][9] .is_wysiwyg = "true";
defparam \openrows[1][9] .power_up = "low";

dffeas \openrows[0][9] (
	.clk(clk),
	.d(\openrows~422_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][9]~q ),
	.prn(vcc));
defparam \openrows[0][9] .is_wysiwyg = "true";
defparam \openrows[0][9] .power_up = "low";

cycloneiii_lcell_comb \Mux3~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][9]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][9]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

dffeas \openrows[3][9] (
	.clk(clk),
	.d(\openrows~422_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][9]~q ),
	.prn(vcc));
defparam \openrows[3][9] .is_wysiwyg = "true";
defparam \openrows[3][9] .power_up = "low";

cycloneiii_lcell_comb \openrows~423 (
	.dataa(row_addr_this_4),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~423_combout ),
	.cout());
defparam \openrows~423 .lut_mask = 16'hAFFF;
defparam \openrows~423 .sum_lutc_input = "datac";

dffeas \openrows[1][4] (
	.clk(clk),
	.d(\openrows~423_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][4]~q ),
	.prn(vcc));
defparam \openrows[1][4] .is_wysiwyg = "true";
defparam \openrows[1][4] .power_up = "low";

dffeas \openrows[2][4] (
	.clk(clk),
	.d(\openrows~423_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][4]~q ),
	.prn(vcc));
defparam \openrows[2][4] .is_wysiwyg = "true";
defparam \openrows[2][4] .power_up = "low";

dffeas \openrows[0][4] (
	.clk(clk),
	.d(\openrows~423_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][4]~q ),
	.prn(vcc));
defparam \openrows[0][4] .is_wysiwyg = "true";
defparam \openrows[0][4] .power_up = "low";

cycloneiii_lcell_comb \Mux8~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][4]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][4]~q ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hFFDE;
defparam \Mux8~0 .sum_lutc_input = "datac";

dffeas \openrows[3][4] (
	.clk(clk),
	.d(\openrows~423_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][4]~q ),
	.prn(vcc));
defparam \openrows[3][4] .is_wysiwyg = "true";
defparam \openrows[3][4] .power_up = "low";

cycloneiii_lcell_comb \openrows~424 (
	.dataa(row_addr_this_10),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~424_combout ),
	.cout());
defparam \openrows~424 .lut_mask = 16'hAFFF;
defparam \openrows~424 .sum_lutc_input = "datac";

dffeas \openrows[1][10] (
	.clk(clk),
	.d(\openrows~424_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][10]~q ),
	.prn(vcc));
defparam \openrows[1][10] .is_wysiwyg = "true";
defparam \openrows[1][10] .power_up = "low";

dffeas \openrows[2][10] (
	.clk(clk),
	.d(\openrows~424_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][10]~q ),
	.prn(vcc));
defparam \openrows[2][10] .is_wysiwyg = "true";
defparam \openrows[2][10] .power_up = "low";

dffeas \openrows[0][10] (
	.clk(clk),
	.d(\openrows~424_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][10]~q ),
	.prn(vcc));
defparam \openrows[0][10] .is_wysiwyg = "true";
defparam \openrows[0][10] .power_up = "low";

cycloneiii_lcell_comb \Mux2~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][10]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][10]~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

dffeas \openrows[3][10] (
	.clk(clk),
	.d(\openrows~424_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][10]~q ),
	.prn(vcc));
defparam \openrows[3][10] .is_wysiwyg = "true";
defparam \openrows[3][10] .power_up = "low";

cycloneiii_lcell_comb \openrows~425 (
	.dataa(row_addr_this_3),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~425_combout ),
	.cout());
defparam \openrows~425 .lut_mask = 16'hAFFF;
defparam \openrows~425 .sum_lutc_input = "datac";

dffeas \openrows[2][3] (
	.clk(clk),
	.d(\openrows~425_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][3]~q ),
	.prn(vcc));
defparam \openrows[2][3] .is_wysiwyg = "true";
defparam \openrows[2][3] .power_up = "low";

dffeas \openrows[1][3] (
	.clk(clk),
	.d(\openrows~425_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][3]~q ),
	.prn(vcc));
defparam \openrows[1][3] .is_wysiwyg = "true";
defparam \openrows[1][3] .power_up = "low";

dffeas \openrows[0][3] (
	.clk(clk),
	.d(\openrows~425_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][3]~q ),
	.prn(vcc));
defparam \openrows[0][3] .is_wysiwyg = "true";
defparam \openrows[0][3] .power_up = "low";

cycloneiii_lcell_comb \Mux9~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][3]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][3]~q ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFFDE;
defparam \Mux9~0 .sum_lutc_input = "datac";

dffeas \openrows[3][3] (
	.clk(clk),
	.d(\openrows~425_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][3]~q ),
	.prn(vcc));
defparam \openrows[3][3] .is_wysiwyg = "true";
defparam \openrows[3][3] .power_up = "low";

cycloneiii_lcell_comb \openrows~426 (
	.dataa(row_addr_this_8),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~426_combout ),
	.cout());
defparam \openrows~426 .lut_mask = 16'hAFFF;
defparam \openrows~426 .sum_lutc_input = "datac";

dffeas \openrows[1][8] (
	.clk(clk),
	.d(\openrows~426_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][8]~q ),
	.prn(vcc));
defparam \openrows[1][8] .is_wysiwyg = "true";
defparam \openrows[1][8] .power_up = "low";

dffeas \openrows[2][8] (
	.clk(clk),
	.d(\openrows~426_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][8]~q ),
	.prn(vcc));
defparam \openrows[2][8] .is_wysiwyg = "true";
defparam \openrows[2][8] .power_up = "low";

dffeas \openrows[0][8] (
	.clk(clk),
	.d(\openrows~426_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][8]~q ),
	.prn(vcc));
defparam \openrows[0][8] .is_wysiwyg = "true";
defparam \openrows[0][8] .power_up = "low";

cycloneiii_lcell_comb \Mux4~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][8]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][8]~q ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hFFDE;
defparam \Mux4~0 .sum_lutc_input = "datac";

dffeas \openrows[3][8] (
	.clk(clk),
	.d(\openrows~426_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][8]~q ),
	.prn(vcc));
defparam \openrows[3][8] .is_wysiwyg = "true";
defparam \openrows[3][8] .power_up = "low";

cycloneiii_lcell_comb \openrows~427 (
	.dataa(row_addr_this_0),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~427_combout ),
	.cout());
defparam \openrows~427 .lut_mask = 16'hAFFF;
defparam \openrows~427 .sum_lutc_input = "datac";

dffeas \openrows[1][0] (
	.clk(clk),
	.d(\openrows~427_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][0]~q ),
	.prn(vcc));
defparam \openrows[1][0] .is_wysiwyg = "true";
defparam \openrows[1][0] .power_up = "low";

dffeas \openrows[2][0] (
	.clk(clk),
	.d(\openrows~427_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][0]~q ),
	.prn(vcc));
defparam \openrows[2][0] .is_wysiwyg = "true";
defparam \openrows[2][0] .power_up = "low";

dffeas \openrows[0][0] (
	.clk(clk),
	.d(\openrows~427_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][0]~q ),
	.prn(vcc));
defparam \openrows[0][0] .is_wysiwyg = "true";
defparam \openrows[0][0] .power_up = "low";

cycloneiii_lcell_comb \Mux12~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][0]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][0]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFFDE;
defparam \Mux12~0 .sum_lutc_input = "datac";

dffeas \openrows[3][0] (
	.clk(clk),
	.d(\openrows~427_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][0]~q ),
	.prn(vcc));
defparam \openrows[3][0] .is_wysiwyg = "true";
defparam \openrows[3][0] .power_up = "low";

cycloneiii_lcell_comb \openrows~428 (
	.dataa(row_addr_this_5),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~428_combout ),
	.cout());
defparam \openrows~428 .lut_mask = 16'hAFFF;
defparam \openrows~428 .sum_lutc_input = "datac";

dffeas \openrows[2][5] (
	.clk(clk),
	.d(\openrows~428_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][5]~q ),
	.prn(vcc));
defparam \openrows[2][5] .is_wysiwyg = "true";
defparam \openrows[2][5] .power_up = "low";

dffeas \openrows[1][5] (
	.clk(clk),
	.d(\openrows~428_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][5]~q ),
	.prn(vcc));
defparam \openrows[1][5] .is_wysiwyg = "true";
defparam \openrows[1][5] .power_up = "low";

dffeas \openrows[0][5] (
	.clk(clk),
	.d(\openrows~428_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][5]~q ),
	.prn(vcc));
defparam \openrows[0][5] .is_wysiwyg = "true";
defparam \openrows[0][5] .power_up = "low";

cycloneiii_lcell_comb \Mux7~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][5]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][5]~q ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hFFDE;
defparam \Mux7~0 .sum_lutc_input = "datac";

dffeas \openrows[3][5] (
	.clk(clk),
	.d(\openrows~428_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][5]~q ),
	.prn(vcc));
defparam \openrows[3][5] .is_wysiwyg = "true";
defparam \openrows[3][5] .power_up = "low";

cycloneiii_lcell_comb \openrows~429 (
	.dataa(row_addr_this_7),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~429_combout ),
	.cout());
defparam \openrows~429 .lut_mask = 16'hAFFF;
defparam \openrows~429 .sum_lutc_input = "datac";

dffeas \openrows[2][7] (
	.clk(clk),
	.d(\openrows~429_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][7]~q ),
	.prn(vcc));
defparam \openrows[2][7] .is_wysiwyg = "true";
defparam \openrows[2][7] .power_up = "low";

dffeas \openrows[1][7] (
	.clk(clk),
	.d(\openrows~429_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][7]~q ),
	.prn(vcc));
defparam \openrows[1][7] .is_wysiwyg = "true";
defparam \openrows[1][7] .power_up = "low";

dffeas \openrows[0][7] (
	.clk(clk),
	.d(\openrows~429_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][7]~q ),
	.prn(vcc));
defparam \openrows[0][7] .is_wysiwyg = "true";
defparam \openrows[0][7] .power_up = "low";

cycloneiii_lcell_comb \Mux5~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][7]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][7]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hFFDE;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \openrows[3][7] (
	.clk(clk),
	.d(\openrows~429_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][7]~q ),
	.prn(vcc));
defparam \openrows[3][7] .is_wysiwyg = "true";
defparam \openrows[3][7] .power_up = "low";

cycloneiii_lcell_comb \openrows~430 (
	.dataa(row_addr_this_6),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~430_combout ),
	.cout());
defparam \openrows~430 .lut_mask = 16'hAFFF;
defparam \openrows~430 .sum_lutc_input = "datac";

dffeas \openrows[1][6] (
	.clk(clk),
	.d(\openrows~430_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][6]~q ),
	.prn(vcc));
defparam \openrows[1][6] .is_wysiwyg = "true";
defparam \openrows[1][6] .power_up = "low";

dffeas \openrows[2][6] (
	.clk(clk),
	.d(\openrows~430_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][6]~q ),
	.prn(vcc));
defparam \openrows[2][6] .is_wysiwyg = "true";
defparam \openrows[2][6] .power_up = "low";

dffeas \openrows[0][6] (
	.clk(clk),
	.d(\openrows~430_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][6]~q ),
	.prn(vcc));
defparam \openrows[0][6] .is_wysiwyg = "true";
defparam \openrows[0][6] .power_up = "low";

cycloneiii_lcell_comb \Mux6~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][6]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][6]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hFFDE;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \openrows[3][6] (
	.clk(clk),
	.d(\openrows~430_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][6]~q ),
	.prn(vcc));
defparam \openrows[3][6] .is_wysiwyg = "true";
defparam \openrows[3][6] .power_up = "low";

cycloneiii_lcell_comb \openrows~431 (
	.dataa(row_addr_this_2),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~431_combout ),
	.cout());
defparam \openrows~431 .lut_mask = 16'hAFFF;
defparam \openrows~431 .sum_lutc_input = "datac";

dffeas \openrows[1][2] (
	.clk(clk),
	.d(\openrows~431_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][2]~q ),
	.prn(vcc));
defparam \openrows[1][2] .is_wysiwyg = "true";
defparam \openrows[1][2] .power_up = "low";

dffeas \openrows[2][2] (
	.clk(clk),
	.d(\openrows~431_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][2]~q ),
	.prn(vcc));
defparam \openrows[2][2] .is_wysiwyg = "true";
defparam \openrows[2][2] .power_up = "low";

dffeas \openrows[0][2] (
	.clk(clk),
	.d(\openrows~431_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][2]~q ),
	.prn(vcc));
defparam \openrows[0][2] .is_wysiwyg = "true";
defparam \openrows[0][2] .power_up = "low";

cycloneiii_lcell_comb \Mux10~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][2]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][2]~q ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hFFDE;
defparam \Mux10~0 .sum_lutc_input = "datac";

dffeas \openrows[3][2] (
	.clk(clk),
	.d(\openrows~431_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][2]~q ),
	.prn(vcc));
defparam \openrows[3][2] .is_wysiwyg = "true";
defparam \openrows[3][2] .power_up = "low";

cycloneiii_lcell_comb \openrows~432 (
	.dataa(row_addr_this_11),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~432_combout ),
	.cout());
defparam \openrows~432 .lut_mask = 16'hAFFF;
defparam \openrows~432 .sum_lutc_input = "datac";

dffeas \openrows[2][11] (
	.clk(clk),
	.d(\openrows~432_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][11]~q ),
	.prn(vcc));
defparam \openrows[2][11] .is_wysiwyg = "true";
defparam \openrows[2][11] .power_up = "low";

dffeas \openrows[1][11] (
	.clk(clk),
	.d(\openrows~432_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][11]~q ),
	.prn(vcc));
defparam \openrows[1][11] .is_wysiwyg = "true";
defparam \openrows[1][11] .power_up = "low";

dffeas \openrows[0][11] (
	.clk(clk),
	.d(\openrows~432_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][11]~q ),
	.prn(vcc));
defparam \openrows[0][11] .is_wysiwyg = "true";
defparam \openrows[0][11] .power_up = "low";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\openrows[1][11]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\openrows[0][11]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas \openrows[3][11] (
	.clk(clk),
	.d(\openrows~432_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][11]~q ),
	.prn(vcc));
defparam \openrows[3][11] .is_wysiwyg = "true";
defparam \openrows[3][11] .power_up = "low";

cycloneiii_lcell_comb \openrows~433 (
	.dataa(row_addr_this_12),
	.datab(gnd),
	.datac(doing_pch_all),
	.datad(doing_pch),
	.cin(gnd),
	.combout(\openrows~433_combout ),
	.cout());
defparam \openrows~433 .lut_mask = 16'hAFFF;
defparam \openrows~433 .sum_lutc_input = "datac";

dffeas \openrows[1][12] (
	.clk(clk),
	.d(\openrows~433_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[1][8]~419_combout ),
	.q(\openrows[1][12]~q ),
	.prn(vcc));
defparam \openrows[1][12] .is_wysiwyg = "true";
defparam \openrows[1][12] .power_up = "low";

dffeas \openrows[2][12] (
	.clk(clk),
	.d(\openrows~433_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[2][11]~418_combout ),
	.q(\openrows[2][12]~q ),
	.prn(vcc));
defparam \openrows[2][12] .is_wysiwyg = "true";
defparam \openrows[2][12] .power_up = "low";

dffeas \openrows[0][12] (
	.clk(clk),
	.d(\openrows~433_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[0][2]~420_combout ),
	.q(\openrows[0][12]~q ),
	.prn(vcc));
defparam \openrows[0][12] .is_wysiwyg = "true";
defparam \openrows[0][12] .power_up = "low";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(row_mux_sel_next_0),
	.datab(\openrows[2][12]~q ),
	.datac(row_mux_sel_next_1),
	.datad(\openrows[0][12]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

dffeas \openrows[3][12] (
	.clk(clk),
	.d(\openrows~433_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\openrows[3][5]~421_combout ),
	.q(\openrows[3][12]~q ),
	.prn(vcc));
defparam \openrows[3][12] .is_wysiwyg = "true";
defparam \openrows[3][12] .power_up = "low";

cycloneiii_lcell_comb \Mux13~0 (
	.dataa(row_mux_sel_next_1),
	.datab(\bank_is_open[1]~q ),
	.datac(row_mux_sel_next_0),
	.datad(\bank_is_open[0]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFFDE;
defparam \Mux13~0 .sum_lutc_input = "datac";

endmodule

module altera_ddr_auk_ddr_hp_input_buf (
	pipefull_3,
	clk,
	seq_ac_add_1t_ac_lat_internal,
	ready,
	reset_n,
	write_req,
	accepted,
	pipefull_0,
	pipe_29_0,
	pipe_28_0,
	pipe_27_0,
	pipe_9_0,
	pipe_8_0,
	pipe_19_0,
	pipe_11_0,
	pipe_14_0,
	pipe_20_0,
	pipe_18_0,
	pipe_13_0,
	pipe_15_0,
	pipe_10_0,
	pipe_16_0,
	pipe_17_0,
	pipe_21_0,
	pipe_12_0,
	pipe_22_0,
	pipe_24_0,
	pipe_25_0,
	pipe_0_0,
	pipe_1_0,
	pipe_2_0,
	pipe_3_0,
	pipe_4_0,
	pipe_5_0,
	pipe_6_0,
	pipe_7_0,
	read_req,
	row_addr,
	bank_addr,
	size,
	col_addr)/* synthesis synthesis_greybox=1 */;
output 	pipefull_3;
input 	clk;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ready;
input 	reset_n;
input 	write_req;
input 	accepted;
output 	pipefull_0;
output 	pipe_29_0;
output 	pipe_28_0;
output 	pipe_27_0;
output 	pipe_9_0;
output 	pipe_8_0;
output 	pipe_19_0;
output 	pipe_11_0;
output 	pipe_14_0;
output 	pipe_20_0;
output 	pipe_18_0;
output 	pipe_13_0;
output 	pipe_15_0;
output 	pipe_10_0;
output 	pipe_16_0;
output 	pipe_17_0;
output 	pipe_21_0;
output 	pipe_12_0;
output 	pipe_22_0;
output 	pipe_24_0;
output 	pipe_25_0;
output 	pipe_0_0;
output 	pipe_1_0;
output 	pipe_2_0;
output 	pipe_3_0;
output 	pipe_4_0;
output 	pipe_5_0;
output 	pipe_6_0;
output 	pipe_7_0;
input 	read_req;
input 	[12:0] row_addr;
input 	[1:0] bank_addr;
input 	[1:0] size;
input 	[7:0] col_addr;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \wr_en~1_combout ;
wire \last_entry_written[10]~q ;
wire \last_entry_written[4]~q ;
wire \Equal0~0_combout ;
wire \last_entry_written[9]~q ;
wire \last_entry_written[1]~q ;
wire \Equal0~1_combout ;
wire \last_entry_written[2]~q ;
wire \last_entry_written[13]~q ;
wire \Equal0~2_combout ;
wire \last_entry_written[0]~q ;
wire \last_entry_written[12]~q ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \last_entry_written[11]~q ;
wire \last_entry_written[5]~q ;
wire \Equal0~5_combout ;
wire \last_entry_written[8]~q ;
wire \last_entry_written[3]~q ;
wire \Equal0~6_combout ;
wire \last_entry_written[7]~q ;
wire \last_entry_written[14]~q ;
wire \Equal0~7_combout ;
wire \last_entry_written[6]~q ;
wire \Equal0~8_combout ;
wire \Equal0~9_combout ;


altera_ddr_auk_ddr_hp_custom_fifo my_fifo(
	.pipefull_3(pipefull_3),
	.clock(clk),
	.ready(ready),
	.aclr(reset_n),
	.data({\Equal0~9_combout ,write_req,read_req,gnd,size[1],size[0],gnd,row_addr[12],row_addr[11],row_addr[10],row_addr[9],row_addr[8],row_addr[7],row_addr[6],row_addr[5],row_addr[4],row_addr[3],row_addr[2],row_addr[1],row_addr[0],bank_addr[1],bank_addr[0],col_addr[7],col_addr[6],col_addr[5],col_addr[4],col_addr[3],col_addr[2],col_addr[1],col_addr[0]}),
	.wr_en(\wr_en~1_combout ),
	.accepted(accepted),
	.pipefull_0(pipefull_0),
	.pipe_29_0(pipe_29_0),
	.pipe_28_0(pipe_28_0),
	.pipe_27_0(pipe_27_0),
	.pipe_9_0(pipe_9_0),
	.pipe_8_0(pipe_8_0),
	.pipe_19_0(pipe_19_0),
	.pipe_11_0(pipe_11_0),
	.pipe_14_0(pipe_14_0),
	.pipe_20_0(pipe_20_0),
	.pipe_18_0(pipe_18_0),
	.pipe_13_0(pipe_13_0),
	.pipe_15_0(pipe_15_0),
	.pipe_10_0(pipe_10_0),
	.pipe_16_0(pipe_16_0),
	.pipe_17_0(pipe_17_0),
	.pipe_21_0(pipe_21_0),
	.pipe_12_0(pipe_12_0),
	.pipe_22_0(pipe_22_0),
	.pipe_24_0(pipe_24_0),
	.pipe_25_0(pipe_25_0),
	.pipe_0_0(pipe_0_0),
	.pipe_1_0(pipe_1_0),
	.pipe_2_0(pipe_2_0),
	.pipe_3_0(pipe_3_0),
	.pipe_4_0(pipe_4_0),
	.pipe_5_0(pipe_5_0),
	.pipe_6_0(pipe_6_0),
	.pipe_7_0(pipe_7_0));

cycloneiii_lcell_comb \wr_en~1 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(read_req),
	.datac(write_req),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\wr_en~1_combout ),
	.cout());
defparam \wr_en~1 .lut_mask = 16'hFEFF;
defparam \wr_en~1 .sum_lutc_input = "datac";

dffeas \last_entry_written[10] (
	.clk(clk),
	.d(row_addr[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[10]~q ),
	.prn(vcc));
defparam \last_entry_written[10] .is_wysiwyg = "true";
defparam \last_entry_written[10] .power_up = "low";

dffeas \last_entry_written[4] (
	.clk(clk),
	.d(row_addr[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[4]~q ),
	.prn(vcc));
defparam \last_entry_written[4] .is_wysiwyg = "true";
defparam \last_entry_written[4] .power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\last_entry_written[10]~q ),
	.datab(\last_entry_written[4]~q ),
	.datac(row_addr[2]),
	.datad(row_addr[8]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

dffeas \last_entry_written[9] (
	.clk(clk),
	.d(row_addr[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[9]~q ),
	.prn(vcc));
defparam \last_entry_written[9] .is_wysiwyg = "true";
defparam \last_entry_written[9] .power_up = "low";

dffeas \last_entry_written[1] (
	.clk(clk),
	.d(bank_addr[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[1]~q ),
	.prn(vcc));
defparam \last_entry_written[1] .is_wysiwyg = "true";
defparam \last_entry_written[1] .power_up = "low";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\last_entry_written[9]~q ),
	.datab(\last_entry_written[1]~q ),
	.datac(bank_addr[1]),
	.datad(row_addr[7]),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

dffeas \last_entry_written[2] (
	.clk(clk),
	.d(row_addr[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[2]~q ),
	.prn(vcc));
defparam \last_entry_written[2] .is_wysiwyg = "true";
defparam \last_entry_written[2] .power_up = "low";

dffeas \last_entry_written[13] (
	.clk(clk),
	.d(row_addr[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[13]~q ),
	.prn(vcc));
defparam \last_entry_written[13] .is_wysiwyg = "true";
defparam \last_entry_written[13] .power_up = "low";

cycloneiii_lcell_comb \Equal0~2 (
	.dataa(\last_entry_written[2]~q ),
	.datab(\last_entry_written[13]~q ),
	.datac(row_addr[11]),
	.datad(row_addr[0]),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h6996;
defparam \Equal0~2 .sum_lutc_input = "datac";

dffeas \last_entry_written[0] (
	.clk(clk),
	.d(bank_addr[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[0]~q ),
	.prn(vcc));
defparam \last_entry_written[0] .is_wysiwyg = "true";
defparam \last_entry_written[0] .power_up = "low";

dffeas \last_entry_written[12] (
	.clk(clk),
	.d(row_addr[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[12]~q ),
	.prn(vcc));
defparam \last_entry_written[12] .is_wysiwyg = "true";
defparam \last_entry_written[12] .power_up = "low";

cycloneiii_lcell_comb \Equal0~3 (
	.dataa(\last_entry_written[0]~q ),
	.datab(\last_entry_written[12]~q ),
	.datac(row_addr[10]),
	.datad(bank_addr[0]),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h6996;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~4 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hFFFE;
defparam \Equal0~4 .sum_lutc_input = "datac";

dffeas \last_entry_written[11] (
	.clk(clk),
	.d(row_addr[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[11]~q ),
	.prn(vcc));
defparam \last_entry_written[11] .is_wysiwyg = "true";
defparam \last_entry_written[11] .power_up = "low";

dffeas \last_entry_written[5] (
	.clk(clk),
	.d(row_addr[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[5]~q ),
	.prn(vcc));
defparam \last_entry_written[5] .is_wysiwyg = "true";
defparam \last_entry_written[5] .power_up = "low";

cycloneiii_lcell_comb \Equal0~5 (
	.dataa(\last_entry_written[11]~q ),
	.datab(\last_entry_written[5]~q ),
	.datac(row_addr[3]),
	.datad(row_addr[9]),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'h6996;
defparam \Equal0~5 .sum_lutc_input = "datac";

dffeas \last_entry_written[8] (
	.clk(clk),
	.d(row_addr[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[8]~q ),
	.prn(vcc));
defparam \last_entry_written[8] .is_wysiwyg = "true";
defparam \last_entry_written[8] .power_up = "low";

dffeas \last_entry_written[3] (
	.clk(clk),
	.d(row_addr[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[3]~q ),
	.prn(vcc));
defparam \last_entry_written[3] .is_wysiwyg = "true";
defparam \last_entry_written[3] .power_up = "low";

cycloneiii_lcell_comb \Equal0~6 (
	.dataa(\last_entry_written[8]~q ),
	.datab(\last_entry_written[3]~q ),
	.datac(row_addr[1]),
	.datad(row_addr[6]),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'h6996;
defparam \Equal0~6 .sum_lutc_input = "datac";

dffeas \last_entry_written[7] (
	.clk(clk),
	.d(row_addr[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[7]~q ),
	.prn(vcc));
defparam \last_entry_written[7] .is_wysiwyg = "true";
defparam \last_entry_written[7] .power_up = "low";

dffeas \last_entry_written[14] (
	.clk(clk),
	.d(row_addr[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[14]~q ),
	.prn(vcc));
defparam \last_entry_written[14] .is_wysiwyg = "true";
defparam \last_entry_written[14] .power_up = "low";

cycloneiii_lcell_comb \Equal0~7 (
	.dataa(\last_entry_written[7]~q ),
	.datab(\last_entry_written[14]~q ),
	.datac(row_addr[12]),
	.datad(row_addr[5]),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'h6996;
defparam \Equal0~7 .sum_lutc_input = "datac";

dffeas \last_entry_written[6] (
	.clk(clk),
	.d(row_addr[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_en~1_combout ),
	.q(\last_entry_written[6]~q ),
	.prn(vcc));
defparam \last_entry_written[6] .is_wysiwyg = "true";
defparam \last_entry_written[6] .power_up = "low";

cycloneiii_lcell_comb \Equal0~8 (
	.dataa(\Equal0~7_combout ),
	.datab(\last_entry_written[6]~q ),
	.datac(row_addr[4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hBEBE;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~9 (
	.dataa(\Equal0~4_combout ),
	.datab(\Equal0~5_combout ),
	.datac(\Equal0~6_combout ),
	.datad(\Equal0~8_combout ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFFFE;
defparam \Equal0~9 .sum_lutc_input = "datac";

endmodule

module altera_ddr_auk_ddr_hp_custom_fifo (
	pipefull_3,
	clock,
	ready,
	aclr,
	data,
	wr_en,
	accepted,
	pipefull_0,
	pipe_29_0,
	pipe_28_0,
	pipe_27_0,
	pipe_9_0,
	pipe_8_0,
	pipe_19_0,
	pipe_11_0,
	pipe_14_0,
	pipe_20_0,
	pipe_18_0,
	pipe_13_0,
	pipe_15_0,
	pipe_10_0,
	pipe_16_0,
	pipe_17_0,
	pipe_21_0,
	pipe_12_0,
	pipe_22_0,
	pipe_24_0,
	pipe_25_0,
	pipe_0_0,
	pipe_1_0,
	pipe_2_0,
	pipe_3_0,
	pipe_4_0,
	pipe_5_0,
	pipe_6_0,
	pipe_7_0)/* synthesis synthesis_greybox=1 */;
output 	pipefull_3;
input 	clock;
input 	ready;
input 	aclr;
input 	[29:0] data;
input 	wr_en;
input 	accepted;
output 	pipefull_0;
output 	pipe_29_0;
output 	pipe_28_0;
output 	pipe_27_0;
output 	pipe_9_0;
output 	pipe_8_0;
output 	pipe_19_0;
output 	pipe_11_0;
output 	pipe_14_0;
output 	pipe_20_0;
output 	pipe_18_0;
output 	pipe_13_0;
output 	pipe_15_0;
output 	pipe_10_0;
output 	pipe_16_0;
output 	pipe_17_0;
output 	pipe_21_0;
output 	pipe_12_0;
output 	pipe_22_0;
output 	pipe_24_0;
output 	pipe_25_0;
output 	pipe_0_0;
output 	pipe_1_0;
output 	pipe_2_0;
output 	pipe_3_0;
output 	pipe_4_0;
output 	pipe_5_0;
output 	pipe_6_0;
output 	pipe_7_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \pipe[2][29]~q ;
wire \pipe[2][28]~q ;
wire \pipe[2][27]~q ;
wire \pipe[2][9]~q ;
wire \pipe[2][8]~q ;
wire \pipe[2][19]~q ;
wire \pipe[2][11]~q ;
wire \pipe[2][14]~q ;
wire \pipe[2][20]~q ;
wire \pipe[2][18]~q ;
wire \pipe[2][13]~q ;
wire \pipe[2][15]~q ;
wire \pipe[2][10]~q ;
wire \pipe[2][16]~q ;
wire \pipe[2][17]~q ;
wire \pipe[2][21]~q ;
wire \pipe[2][12]~q ;
wire \pipe[2][22]~q ;
wire \pipe[3][29]~q ;
wire \pipe~128_combout ;
wire \process_2~0_combout ;
wire \pipe[3][28]~q ;
wire \pipe~129_combout ;
wire \pipe[2][24]~q ;
wire \pipe[2][25]~q ;
wire \pipe[3][27]~q ;
wire \pipe~132_combout ;
wire \pipe[3][9]~q ;
wire \pipe~141_combout ;
wire \pipe[3][8]~q ;
wire \pipe~142_combout ;
wire \pipe[3][19]~q ;
wire \pipe~143_combout ;
wire \pipe[3][11]~q ;
wire \pipe~144_combout ;
wire \pipe[3][14]~q ;
wire \pipe~145_combout ;
wire \pipe[3][20]~q ;
wire \pipe~146_combout ;
wire \pipe[3][18]~q ;
wire \pipe~147_combout ;
wire \pipe[3][13]~q ;
wire \pipe~148_combout ;
wire \pipe[3][15]~q ;
wire \pipe~149_combout ;
wire \pipe[3][10]~q ;
wire \pipe~150_combout ;
wire \pipe[3][16]~q ;
wire \pipe~151_combout ;
wire \pipe[3][17]~q ;
wire \pipe~152_combout ;
wire \pipe[3][21]~q ;
wire \pipe~153_combout ;
wire \pipe[3][12]~q ;
wire \pipe~154_combout ;
wire \pipe[3][22]~q ;
wire \pipe~155_combout ;
wire \process_0~1_combout ;
wire \pipe[3][24]~q ;
wire \pipe~156_combout ;
wire \pipe[3][25]~q ;
wire \pipe~157_combout ;
wire \pipe[2][0]~q ;
wire \pipe[2][1]~q ;
wire \pipe[2][2]~q ;
wire \pipe[2][3]~q ;
wire \pipe[2][4]~q ;
wire \pipe[2][5]~q ;
wire \pipe[2][6]~q ;
wire \pipe[2][7]~q ;
wire \pipe[3][0]~q ;
wire \pipe~166_combout ;
wire \pipe[3][1]~q ;
wire \pipe~167_combout ;
wire \pipe[3][2]~q ;
wire \pipe~168_combout ;
wire \pipe[3][3]~q ;
wire \pipe~169_combout ;
wire \pipe[3][4]~q ;
wire \pipe~170_combout ;
wire \pipe[3][5]~q ;
wire \pipe~171_combout ;
wire \pipe[3][6]~q ;
wire \pipe~172_combout ;
wire \pipe[3][7]~q ;
wire \pipe~173_combout ;
wire \pipefull~11_combout ;
wire \process_0~2_combout ;
wire \pipefull[1]~q ;
wire \pipefull~10_combout ;
wire \pipefull[2]~q ;
wire \pipefull[3]~9_combout ;
wire \pipefull[0]~12_combout ;
wire \pipe~108_combout ;
wire \process_1~0_combout ;
wire \pipe[1][29]~q ;
wire \pipe~90_combout ;
wire \process_0~0_combout ;
wire \pipe~109_combout ;
wire \pipe[1][28]~q ;
wire \pipe~91_combout ;
wire \pipe~112_combout ;
wire \pipe[1][27]~q ;
wire \pipe~92_combout ;
wire \pipe~113_combout ;
wire \pipe[1][9]~q ;
wire \pipe~93_combout ;
wire \pipe~114_combout ;
wire \pipe[1][8]~q ;
wire \pipe~94_combout ;
wire \pipe~115_combout ;
wire \pipe[1][19]~q ;
wire \pipe~95_combout ;
wire \pipe~116_combout ;
wire \pipe[1][11]~q ;
wire \pipe~96_combout ;
wire \pipe~117_combout ;
wire \pipe[1][14]~q ;
wire \pipe~97_combout ;
wire \pipe~118_combout ;
wire \pipe[1][20]~q ;
wire \pipe~98_combout ;
wire \pipe~119_combout ;
wire \pipe[1][18]~q ;
wire \pipe~99_combout ;
wire \pipe~120_combout ;
wire \pipe[1][13]~q ;
wire \pipe~100_combout ;
wire \pipe~121_combout ;
wire \pipe[1][15]~q ;
wire \pipe~101_combout ;
wire \pipe~122_combout ;
wire \pipe[1][10]~q ;
wire \pipe~102_combout ;
wire \pipe~123_combout ;
wire \pipe[1][16]~q ;
wire \pipe~103_combout ;
wire \pipe~124_combout ;
wire \pipe[1][17]~q ;
wire \pipe~104_combout ;
wire \pipe~125_combout ;
wire \pipe[1][21]~q ;
wire \pipe~105_combout ;
wire \pipe~126_combout ;
wire \pipe[1][12]~q ;
wire \pipe~106_combout ;
wire \pipe~127_combout ;
wire \pipe[1][22]~q ;
wire \pipe~107_combout ;
wire \pipe~130_combout ;
wire \pipe[1][24]~q ;
wire \pipe~110_combout ;
wire \pipe~131_combout ;
wire \pipe[1][25]~q ;
wire \pipe~111_combout ;
wire \pipe~158_combout ;
wire \pipe[1][0]~q ;
wire \pipe~133_combout ;
wire \pipe~159_combout ;
wire \pipe[1][1]~q ;
wire \pipe~134_combout ;
wire \pipe~160_combout ;
wire \pipe[1][2]~q ;
wire \pipe~135_combout ;
wire \pipe~161_combout ;
wire \pipe[1][3]~q ;
wire \pipe~136_combout ;
wire \pipe~162_combout ;
wire \pipe[1][4]~q ;
wire \pipe~137_combout ;
wire \pipe~163_combout ;
wire \pipe[1][5]~q ;
wire \pipe~138_combout ;
wire \pipe~164_combout ;
wire \pipe[1][6]~q ;
wire \pipe~139_combout ;
wire \pipe~165_combout ;
wire \pipe[1][7]~q ;
wire \pipe~140_combout ;


dffeas \pipe[2][29] (
	.clk(clock),
	.d(\pipe~128_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][29]~q ),
	.prn(vcc));
defparam \pipe[2][29] .is_wysiwyg = "true";
defparam \pipe[2][29] .power_up = "low";

dffeas \pipe[2][28] (
	.clk(clock),
	.d(\pipe~129_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][28]~q ),
	.prn(vcc));
defparam \pipe[2][28] .is_wysiwyg = "true";
defparam \pipe[2][28] .power_up = "low";

dffeas \pipe[2][27] (
	.clk(clock),
	.d(\pipe~132_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][27]~q ),
	.prn(vcc));
defparam \pipe[2][27] .is_wysiwyg = "true";
defparam \pipe[2][27] .power_up = "low";

dffeas \pipe[2][9] (
	.clk(clock),
	.d(\pipe~141_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][9]~q ),
	.prn(vcc));
defparam \pipe[2][9] .is_wysiwyg = "true";
defparam \pipe[2][9] .power_up = "low";

dffeas \pipe[2][8] (
	.clk(clock),
	.d(\pipe~142_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][8]~q ),
	.prn(vcc));
defparam \pipe[2][8] .is_wysiwyg = "true";
defparam \pipe[2][8] .power_up = "low";

dffeas \pipe[2][19] (
	.clk(clock),
	.d(\pipe~143_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][19]~q ),
	.prn(vcc));
defparam \pipe[2][19] .is_wysiwyg = "true";
defparam \pipe[2][19] .power_up = "low";

dffeas \pipe[2][11] (
	.clk(clock),
	.d(\pipe~144_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][11]~q ),
	.prn(vcc));
defparam \pipe[2][11] .is_wysiwyg = "true";
defparam \pipe[2][11] .power_up = "low";

dffeas \pipe[2][14] (
	.clk(clock),
	.d(\pipe~145_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][14]~q ),
	.prn(vcc));
defparam \pipe[2][14] .is_wysiwyg = "true";
defparam \pipe[2][14] .power_up = "low";

dffeas \pipe[2][20] (
	.clk(clock),
	.d(\pipe~146_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][20]~q ),
	.prn(vcc));
defparam \pipe[2][20] .is_wysiwyg = "true";
defparam \pipe[2][20] .power_up = "low";

dffeas \pipe[2][18] (
	.clk(clock),
	.d(\pipe~147_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][18]~q ),
	.prn(vcc));
defparam \pipe[2][18] .is_wysiwyg = "true";
defparam \pipe[2][18] .power_up = "low";

dffeas \pipe[2][13] (
	.clk(clock),
	.d(\pipe~148_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][13]~q ),
	.prn(vcc));
defparam \pipe[2][13] .is_wysiwyg = "true";
defparam \pipe[2][13] .power_up = "low";

dffeas \pipe[2][15] (
	.clk(clock),
	.d(\pipe~149_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][15]~q ),
	.prn(vcc));
defparam \pipe[2][15] .is_wysiwyg = "true";
defparam \pipe[2][15] .power_up = "low";

dffeas \pipe[2][10] (
	.clk(clock),
	.d(\pipe~150_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][10]~q ),
	.prn(vcc));
defparam \pipe[2][10] .is_wysiwyg = "true";
defparam \pipe[2][10] .power_up = "low";

dffeas \pipe[2][16] (
	.clk(clock),
	.d(\pipe~151_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][16]~q ),
	.prn(vcc));
defparam \pipe[2][16] .is_wysiwyg = "true";
defparam \pipe[2][16] .power_up = "low";

dffeas \pipe[2][17] (
	.clk(clock),
	.d(\pipe~152_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][17]~q ),
	.prn(vcc));
defparam \pipe[2][17] .is_wysiwyg = "true";
defparam \pipe[2][17] .power_up = "low";

dffeas \pipe[2][21] (
	.clk(clock),
	.d(\pipe~153_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][21]~q ),
	.prn(vcc));
defparam \pipe[2][21] .is_wysiwyg = "true";
defparam \pipe[2][21] .power_up = "low";

dffeas \pipe[2][12] (
	.clk(clock),
	.d(\pipe~154_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][12]~q ),
	.prn(vcc));
defparam \pipe[2][12] .is_wysiwyg = "true";
defparam \pipe[2][12] .power_up = "low";

dffeas \pipe[2][22] (
	.clk(clock),
	.d(\pipe~155_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][22]~q ),
	.prn(vcc));
defparam \pipe[2][22] .is_wysiwyg = "true";
defparam \pipe[2][22] .power_up = "low";

dffeas \pipe[3][29] (
	.clk(clock),
	.d(data[29]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][29]~q ),
	.prn(vcc));
defparam \pipe[3][29] .is_wysiwyg = "true";
defparam \pipe[3][29] .power_up = "low";

cycloneiii_lcell_comb \pipe~128 (
	.dataa(\pipe[3][29]~q ),
	.datab(data[29]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~128_combout ),
	.cout());
defparam \pipe~128 .lut_mask = 16'hAACC;
defparam \pipe~128 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_2~0 (
	.dataa(accepted),
	.datab(gnd),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\process_2~0_combout ),
	.cout());
defparam \process_2~0 .lut_mask = 16'hAAFF;
defparam \process_2~0 .sum_lutc_input = "datac";

dffeas \pipe[3][28] (
	.clk(clock),
	.d(data[28]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][28]~q ),
	.prn(vcc));
defparam \pipe[3][28] .is_wysiwyg = "true";
defparam \pipe[3][28] .power_up = "low";

cycloneiii_lcell_comb \pipe~129 (
	.dataa(\pipe[3][28]~q ),
	.datab(data[28]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~129_combout ),
	.cout());
defparam \pipe~129 .lut_mask = 16'hAACC;
defparam \pipe~129 .sum_lutc_input = "datac";

dffeas \pipe[2][24] (
	.clk(clock),
	.d(\pipe~156_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][24]~q ),
	.prn(vcc));
defparam \pipe[2][24] .is_wysiwyg = "true";
defparam \pipe[2][24] .power_up = "low";

dffeas \pipe[2][25] (
	.clk(clock),
	.d(\pipe~157_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][25]~q ),
	.prn(vcc));
defparam \pipe[2][25] .is_wysiwyg = "true";
defparam \pipe[2][25] .power_up = "low";

dffeas \pipe[3][27] (
	.clk(clock),
	.d(data[27]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][27]~q ),
	.prn(vcc));
defparam \pipe[3][27] .is_wysiwyg = "true";
defparam \pipe[3][27] .power_up = "low";

cycloneiii_lcell_comb \pipe~132 (
	.dataa(\pipe[3][27]~q ),
	.datab(data[27]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~132_combout ),
	.cout());
defparam \pipe~132 .lut_mask = 16'hAACC;
defparam \pipe~132 .sum_lutc_input = "datac";

dffeas \pipe[3][9] (
	.clk(clock),
	.d(data[9]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][9]~q ),
	.prn(vcc));
defparam \pipe[3][9] .is_wysiwyg = "true";
defparam \pipe[3][9] .power_up = "low";

cycloneiii_lcell_comb \pipe~141 (
	.dataa(\pipe[3][9]~q ),
	.datab(data[9]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~141_combout ),
	.cout());
defparam \pipe~141 .lut_mask = 16'hAACC;
defparam \pipe~141 .sum_lutc_input = "datac";

dffeas \pipe[3][8] (
	.clk(clock),
	.d(data[8]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][8]~q ),
	.prn(vcc));
defparam \pipe[3][8] .is_wysiwyg = "true";
defparam \pipe[3][8] .power_up = "low";

cycloneiii_lcell_comb \pipe~142 (
	.dataa(\pipe[3][8]~q ),
	.datab(data[8]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~142_combout ),
	.cout());
defparam \pipe~142 .lut_mask = 16'hAACC;
defparam \pipe~142 .sum_lutc_input = "datac";

dffeas \pipe[3][19] (
	.clk(clock),
	.d(data[19]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][19]~q ),
	.prn(vcc));
defparam \pipe[3][19] .is_wysiwyg = "true";
defparam \pipe[3][19] .power_up = "low";

cycloneiii_lcell_comb \pipe~143 (
	.dataa(\pipe[3][19]~q ),
	.datab(data[19]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~143_combout ),
	.cout());
defparam \pipe~143 .lut_mask = 16'hAACC;
defparam \pipe~143 .sum_lutc_input = "datac";

dffeas \pipe[3][11] (
	.clk(clock),
	.d(data[11]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][11]~q ),
	.prn(vcc));
defparam \pipe[3][11] .is_wysiwyg = "true";
defparam \pipe[3][11] .power_up = "low";

cycloneiii_lcell_comb \pipe~144 (
	.dataa(\pipe[3][11]~q ),
	.datab(data[11]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~144_combout ),
	.cout());
defparam \pipe~144 .lut_mask = 16'hAACC;
defparam \pipe~144 .sum_lutc_input = "datac";

dffeas \pipe[3][14] (
	.clk(clock),
	.d(data[14]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][14]~q ),
	.prn(vcc));
defparam \pipe[3][14] .is_wysiwyg = "true";
defparam \pipe[3][14] .power_up = "low";

cycloneiii_lcell_comb \pipe~145 (
	.dataa(\pipe[3][14]~q ),
	.datab(data[14]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~145_combout ),
	.cout());
defparam \pipe~145 .lut_mask = 16'hAACC;
defparam \pipe~145 .sum_lutc_input = "datac";

dffeas \pipe[3][20] (
	.clk(clock),
	.d(data[20]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][20]~q ),
	.prn(vcc));
defparam \pipe[3][20] .is_wysiwyg = "true";
defparam \pipe[3][20] .power_up = "low";

cycloneiii_lcell_comb \pipe~146 (
	.dataa(\pipe[3][20]~q ),
	.datab(data[20]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~146_combout ),
	.cout());
defparam \pipe~146 .lut_mask = 16'hAACC;
defparam \pipe~146 .sum_lutc_input = "datac";

dffeas \pipe[3][18] (
	.clk(clock),
	.d(data[18]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][18]~q ),
	.prn(vcc));
defparam \pipe[3][18] .is_wysiwyg = "true";
defparam \pipe[3][18] .power_up = "low";

cycloneiii_lcell_comb \pipe~147 (
	.dataa(\pipe[3][18]~q ),
	.datab(data[18]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~147_combout ),
	.cout());
defparam \pipe~147 .lut_mask = 16'hAACC;
defparam \pipe~147 .sum_lutc_input = "datac";

dffeas \pipe[3][13] (
	.clk(clock),
	.d(data[13]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][13]~q ),
	.prn(vcc));
defparam \pipe[3][13] .is_wysiwyg = "true";
defparam \pipe[3][13] .power_up = "low";

cycloneiii_lcell_comb \pipe~148 (
	.dataa(\pipe[3][13]~q ),
	.datab(data[13]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~148_combout ),
	.cout());
defparam \pipe~148 .lut_mask = 16'hAACC;
defparam \pipe~148 .sum_lutc_input = "datac";

dffeas \pipe[3][15] (
	.clk(clock),
	.d(data[15]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][15]~q ),
	.prn(vcc));
defparam \pipe[3][15] .is_wysiwyg = "true";
defparam \pipe[3][15] .power_up = "low";

cycloneiii_lcell_comb \pipe~149 (
	.dataa(\pipe[3][15]~q ),
	.datab(data[15]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~149_combout ),
	.cout());
defparam \pipe~149 .lut_mask = 16'hAACC;
defparam \pipe~149 .sum_lutc_input = "datac";

dffeas \pipe[3][10] (
	.clk(clock),
	.d(data[10]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][10]~q ),
	.prn(vcc));
defparam \pipe[3][10] .is_wysiwyg = "true";
defparam \pipe[3][10] .power_up = "low";

cycloneiii_lcell_comb \pipe~150 (
	.dataa(\pipe[3][10]~q ),
	.datab(data[10]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~150_combout ),
	.cout());
defparam \pipe~150 .lut_mask = 16'hAACC;
defparam \pipe~150 .sum_lutc_input = "datac";

dffeas \pipe[3][16] (
	.clk(clock),
	.d(data[16]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][16]~q ),
	.prn(vcc));
defparam \pipe[3][16] .is_wysiwyg = "true";
defparam \pipe[3][16] .power_up = "low";

cycloneiii_lcell_comb \pipe~151 (
	.dataa(\pipe[3][16]~q ),
	.datab(data[16]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~151_combout ),
	.cout());
defparam \pipe~151 .lut_mask = 16'hAACC;
defparam \pipe~151 .sum_lutc_input = "datac";

dffeas \pipe[3][17] (
	.clk(clock),
	.d(data[17]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][17]~q ),
	.prn(vcc));
defparam \pipe[3][17] .is_wysiwyg = "true";
defparam \pipe[3][17] .power_up = "low";

cycloneiii_lcell_comb \pipe~152 (
	.dataa(\pipe[3][17]~q ),
	.datab(data[17]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~152_combout ),
	.cout());
defparam \pipe~152 .lut_mask = 16'hAACC;
defparam \pipe~152 .sum_lutc_input = "datac";

dffeas \pipe[3][21] (
	.clk(clock),
	.d(data[21]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][21]~q ),
	.prn(vcc));
defparam \pipe[3][21] .is_wysiwyg = "true";
defparam \pipe[3][21] .power_up = "low";

cycloneiii_lcell_comb \pipe~153 (
	.dataa(\pipe[3][21]~q ),
	.datab(data[21]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~153_combout ),
	.cout());
defparam \pipe~153 .lut_mask = 16'hAACC;
defparam \pipe~153 .sum_lutc_input = "datac";

dffeas \pipe[3][12] (
	.clk(clock),
	.d(data[12]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][12]~q ),
	.prn(vcc));
defparam \pipe[3][12] .is_wysiwyg = "true";
defparam \pipe[3][12] .power_up = "low";

cycloneiii_lcell_comb \pipe~154 (
	.dataa(\pipe[3][12]~q ),
	.datab(data[12]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~154_combout ),
	.cout());
defparam \pipe~154 .lut_mask = 16'hAACC;
defparam \pipe~154 .sum_lutc_input = "datac";

dffeas \pipe[3][22] (
	.clk(clock),
	.d(data[22]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][22]~q ),
	.prn(vcc));
defparam \pipe[3][22] .is_wysiwyg = "true";
defparam \pipe[3][22] .power_up = "low";

cycloneiii_lcell_comb \pipe~155 (
	.dataa(\pipe[3][22]~q ),
	.datab(data[22]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~155_combout ),
	.cout());
defparam \pipe~155 .lut_mask = 16'hAACC;
defparam \pipe~155 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_0~1 (
	.dataa(accepted),
	.datab(gnd),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
defparam \process_0~1 .lut_mask = 16'hAAFF;
defparam \process_0~1 .sum_lutc_input = "datac";

dffeas \pipe[3][24] (
	.clk(clock),
	.d(data[24]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][24]~q ),
	.prn(vcc));
defparam \pipe[3][24] .is_wysiwyg = "true";
defparam \pipe[3][24] .power_up = "low";

cycloneiii_lcell_comb \pipe~156 (
	.dataa(\pipe[3][24]~q ),
	.datab(data[24]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~156_combout ),
	.cout());
defparam \pipe~156 .lut_mask = 16'hAACC;
defparam \pipe~156 .sum_lutc_input = "datac";

dffeas \pipe[3][25] (
	.clk(clock),
	.d(data[25]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][25]~q ),
	.prn(vcc));
defparam \pipe[3][25] .is_wysiwyg = "true";
defparam \pipe[3][25] .power_up = "low";

cycloneiii_lcell_comb \pipe~157 (
	.dataa(\pipe[3][25]~q ),
	.datab(data[25]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~157_combout ),
	.cout());
defparam \pipe~157 .lut_mask = 16'hAACC;
defparam \pipe~157 .sum_lutc_input = "datac";

dffeas \pipe[2][0] (
	.clk(clock),
	.d(\pipe~166_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][0]~q ),
	.prn(vcc));
defparam \pipe[2][0] .is_wysiwyg = "true";
defparam \pipe[2][0] .power_up = "low";

dffeas \pipe[2][1] (
	.clk(clock),
	.d(\pipe~167_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][1]~q ),
	.prn(vcc));
defparam \pipe[2][1] .is_wysiwyg = "true";
defparam \pipe[2][1] .power_up = "low";

dffeas \pipe[2][2] (
	.clk(clock),
	.d(\pipe~168_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][2]~q ),
	.prn(vcc));
defparam \pipe[2][2] .is_wysiwyg = "true";
defparam \pipe[2][2] .power_up = "low";

dffeas \pipe[2][3] (
	.clk(clock),
	.d(\pipe~169_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][3]~q ),
	.prn(vcc));
defparam \pipe[2][3] .is_wysiwyg = "true";
defparam \pipe[2][3] .power_up = "low";

dffeas \pipe[2][4] (
	.clk(clock),
	.d(\pipe~170_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][4]~q ),
	.prn(vcc));
defparam \pipe[2][4] .is_wysiwyg = "true";
defparam \pipe[2][4] .power_up = "low";

dffeas \pipe[2][5] (
	.clk(clock),
	.d(\pipe~171_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][5]~q ),
	.prn(vcc));
defparam \pipe[2][5] .is_wysiwyg = "true";
defparam \pipe[2][5] .power_up = "low";

dffeas \pipe[2][6] (
	.clk(clock),
	.d(\pipe~172_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][6]~q ),
	.prn(vcc));
defparam \pipe[2][6] .is_wysiwyg = "true";
defparam \pipe[2][6] .power_up = "low";

dffeas \pipe[2][7] (
	.clk(clock),
	.d(\pipe~173_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_2~0_combout ),
	.q(\pipe[2][7]~q ),
	.prn(vcc));
defparam \pipe[2][7] .is_wysiwyg = "true";
defparam \pipe[2][7] .power_up = "low";

dffeas \pipe[3][0] (
	.clk(clock),
	.d(data[0]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][0]~q ),
	.prn(vcc));
defparam \pipe[3][0] .is_wysiwyg = "true";
defparam \pipe[3][0] .power_up = "low";

cycloneiii_lcell_comb \pipe~166 (
	.dataa(\pipe[3][0]~q ),
	.datab(data[0]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~166_combout ),
	.cout());
defparam \pipe~166 .lut_mask = 16'hAACC;
defparam \pipe~166 .sum_lutc_input = "datac";

dffeas \pipe[3][1] (
	.clk(clock),
	.d(data[1]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][1]~q ),
	.prn(vcc));
defparam \pipe[3][1] .is_wysiwyg = "true";
defparam \pipe[3][1] .power_up = "low";

cycloneiii_lcell_comb \pipe~167 (
	.dataa(\pipe[3][1]~q ),
	.datab(data[1]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~167_combout ),
	.cout());
defparam \pipe~167 .lut_mask = 16'hAACC;
defparam \pipe~167 .sum_lutc_input = "datac";

dffeas \pipe[3][2] (
	.clk(clock),
	.d(data[2]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][2]~q ),
	.prn(vcc));
defparam \pipe[3][2] .is_wysiwyg = "true";
defparam \pipe[3][2] .power_up = "low";

cycloneiii_lcell_comb \pipe~168 (
	.dataa(\pipe[3][2]~q ),
	.datab(data[2]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~168_combout ),
	.cout());
defparam \pipe~168 .lut_mask = 16'hAACC;
defparam \pipe~168 .sum_lutc_input = "datac";

dffeas \pipe[3][3] (
	.clk(clock),
	.d(data[3]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][3]~q ),
	.prn(vcc));
defparam \pipe[3][3] .is_wysiwyg = "true";
defparam \pipe[3][3] .power_up = "low";

cycloneiii_lcell_comb \pipe~169 (
	.dataa(\pipe[3][3]~q ),
	.datab(data[3]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~169_combout ),
	.cout());
defparam \pipe~169 .lut_mask = 16'hAACC;
defparam \pipe~169 .sum_lutc_input = "datac";

dffeas \pipe[3][4] (
	.clk(clock),
	.d(data[4]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][4]~q ),
	.prn(vcc));
defparam \pipe[3][4] .is_wysiwyg = "true";
defparam \pipe[3][4] .power_up = "low";

cycloneiii_lcell_comb \pipe~170 (
	.dataa(\pipe[3][4]~q ),
	.datab(data[4]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~170_combout ),
	.cout());
defparam \pipe~170 .lut_mask = 16'hAACC;
defparam \pipe~170 .sum_lutc_input = "datac";

dffeas \pipe[3][5] (
	.clk(clock),
	.d(data[5]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][5]~q ),
	.prn(vcc));
defparam \pipe[3][5] .is_wysiwyg = "true";
defparam \pipe[3][5] .power_up = "low";

cycloneiii_lcell_comb \pipe~171 (
	.dataa(\pipe[3][5]~q ),
	.datab(data[5]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~171_combout ),
	.cout());
defparam \pipe~171 .lut_mask = 16'hAACC;
defparam \pipe~171 .sum_lutc_input = "datac";

dffeas \pipe[3][6] (
	.clk(clock),
	.d(data[6]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][6]~q ),
	.prn(vcc));
defparam \pipe[3][6] .is_wysiwyg = "true";
defparam \pipe[3][6] .power_up = "low";

cycloneiii_lcell_comb \pipe~172 (
	.dataa(\pipe[3][6]~q ),
	.datab(data[6]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~172_combout ),
	.cout());
defparam \pipe~172 .lut_mask = 16'hAACC;
defparam \pipe~172 .sum_lutc_input = "datac";

dffeas \pipe[3][7] (
	.clk(clock),
	.d(data[7]),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.q(\pipe[3][7]~q ),
	.prn(vcc));
defparam \pipe[3][7] .is_wysiwyg = "true";
defparam \pipe[3][7] .power_up = "low";

cycloneiii_lcell_comb \pipe~173 (
	.dataa(\pipe[3][7]~q ),
	.datab(data[7]),
	.datac(gnd),
	.datad(pipefull_3),
	.cin(gnd),
	.combout(\pipe~173_combout ),
	.cout());
defparam \pipe~173 .lut_mask = 16'hAACC;
defparam \pipe~173 .sum_lutc_input = "datac";

dffeas \pipefull[3] (
	.clk(clock),
	.d(\pipefull[3]~9_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(accepted),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_3),
	.prn(vcc));
defparam \pipefull[3] .is_wysiwyg = "true";
defparam \pipefull[3] .power_up = "low";

dffeas \pipefull[0] (
	.clk(clock),
	.d(\pipefull[0]~12_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_0),
	.prn(vcc));
defparam \pipefull[0] .is_wysiwyg = "true";
defparam \pipefull[0] .power_up = "low";

dffeas \pipe[0][29] (
	.clk(clock),
	.d(\pipe~90_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_29_0),
	.prn(vcc));
defparam \pipe[0][29] .is_wysiwyg = "true";
defparam \pipe[0][29] .power_up = "low";

dffeas \pipe[0][28] (
	.clk(clock),
	.d(\pipe~91_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_28_0),
	.prn(vcc));
defparam \pipe[0][28] .is_wysiwyg = "true";
defparam \pipe[0][28] .power_up = "low";

dffeas \pipe[0][27] (
	.clk(clock),
	.d(\pipe~92_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_27_0),
	.prn(vcc));
defparam \pipe[0][27] .is_wysiwyg = "true";
defparam \pipe[0][27] .power_up = "low";

dffeas \pipe[0][9] (
	.clk(clock),
	.d(\pipe~93_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_9_0),
	.prn(vcc));
defparam \pipe[0][9] .is_wysiwyg = "true";
defparam \pipe[0][9] .power_up = "low";

dffeas \pipe[0][8] (
	.clk(clock),
	.d(\pipe~94_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_8_0),
	.prn(vcc));
defparam \pipe[0][8] .is_wysiwyg = "true";
defparam \pipe[0][8] .power_up = "low";

dffeas \pipe[0][19] (
	.clk(clock),
	.d(\pipe~95_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_19_0),
	.prn(vcc));
defparam \pipe[0][19] .is_wysiwyg = "true";
defparam \pipe[0][19] .power_up = "low";

dffeas \pipe[0][11] (
	.clk(clock),
	.d(\pipe~96_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_11_0),
	.prn(vcc));
defparam \pipe[0][11] .is_wysiwyg = "true";
defparam \pipe[0][11] .power_up = "low";

dffeas \pipe[0][14] (
	.clk(clock),
	.d(\pipe~97_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_14_0),
	.prn(vcc));
defparam \pipe[0][14] .is_wysiwyg = "true";
defparam \pipe[0][14] .power_up = "low";

dffeas \pipe[0][20] (
	.clk(clock),
	.d(\pipe~98_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_20_0),
	.prn(vcc));
defparam \pipe[0][20] .is_wysiwyg = "true";
defparam \pipe[0][20] .power_up = "low";

dffeas \pipe[0][18] (
	.clk(clock),
	.d(\pipe~99_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_18_0),
	.prn(vcc));
defparam \pipe[0][18] .is_wysiwyg = "true";
defparam \pipe[0][18] .power_up = "low";

dffeas \pipe[0][13] (
	.clk(clock),
	.d(\pipe~100_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_13_0),
	.prn(vcc));
defparam \pipe[0][13] .is_wysiwyg = "true";
defparam \pipe[0][13] .power_up = "low";

dffeas \pipe[0][15] (
	.clk(clock),
	.d(\pipe~101_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_15_0),
	.prn(vcc));
defparam \pipe[0][15] .is_wysiwyg = "true";
defparam \pipe[0][15] .power_up = "low";

dffeas \pipe[0][10] (
	.clk(clock),
	.d(\pipe~102_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_10_0),
	.prn(vcc));
defparam \pipe[0][10] .is_wysiwyg = "true";
defparam \pipe[0][10] .power_up = "low";

dffeas \pipe[0][16] (
	.clk(clock),
	.d(\pipe~103_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_16_0),
	.prn(vcc));
defparam \pipe[0][16] .is_wysiwyg = "true";
defparam \pipe[0][16] .power_up = "low";

dffeas \pipe[0][17] (
	.clk(clock),
	.d(\pipe~104_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_17_0),
	.prn(vcc));
defparam \pipe[0][17] .is_wysiwyg = "true";
defparam \pipe[0][17] .power_up = "low";

dffeas \pipe[0][21] (
	.clk(clock),
	.d(\pipe~105_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_21_0),
	.prn(vcc));
defparam \pipe[0][21] .is_wysiwyg = "true";
defparam \pipe[0][21] .power_up = "low";

dffeas \pipe[0][12] (
	.clk(clock),
	.d(\pipe~106_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_12_0),
	.prn(vcc));
defparam \pipe[0][12] .is_wysiwyg = "true";
defparam \pipe[0][12] .power_up = "low";

dffeas \pipe[0][22] (
	.clk(clock),
	.d(\pipe~107_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_22_0),
	.prn(vcc));
defparam \pipe[0][22] .is_wysiwyg = "true";
defparam \pipe[0][22] .power_up = "low";

dffeas \pipe[0][24] (
	.clk(clock),
	.d(\pipe~110_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_24_0),
	.prn(vcc));
defparam \pipe[0][24] .is_wysiwyg = "true";
defparam \pipe[0][24] .power_up = "low";

dffeas \pipe[0][25] (
	.clk(clock),
	.d(\pipe~111_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_25_0),
	.prn(vcc));
defparam \pipe[0][25] .is_wysiwyg = "true";
defparam \pipe[0][25] .power_up = "low";

dffeas \pipe[0][0] (
	.clk(clock),
	.d(\pipe~133_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_0_0),
	.prn(vcc));
defparam \pipe[0][0] .is_wysiwyg = "true";
defparam \pipe[0][0] .power_up = "low";

dffeas \pipe[0][1] (
	.clk(clock),
	.d(\pipe~134_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_1_0),
	.prn(vcc));
defparam \pipe[0][1] .is_wysiwyg = "true";
defparam \pipe[0][1] .power_up = "low";

dffeas \pipe[0][2] (
	.clk(clock),
	.d(\pipe~135_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_2_0),
	.prn(vcc));
defparam \pipe[0][2] .is_wysiwyg = "true";
defparam \pipe[0][2] .power_up = "low";

dffeas \pipe[0][3] (
	.clk(clock),
	.d(\pipe~136_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_3_0),
	.prn(vcc));
defparam \pipe[0][3] .is_wysiwyg = "true";
defparam \pipe[0][3] .power_up = "low";

dffeas \pipe[0][4] (
	.clk(clock),
	.d(\pipe~137_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_4_0),
	.prn(vcc));
defparam \pipe[0][4] .is_wysiwyg = "true";
defparam \pipe[0][4] .power_up = "low";

dffeas \pipe[0][5] (
	.clk(clock),
	.d(\pipe~138_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_5_0),
	.prn(vcc));
defparam \pipe[0][5] .is_wysiwyg = "true";
defparam \pipe[0][5] .power_up = "low";

dffeas \pipe[0][6] (
	.clk(clock),
	.d(\pipe~139_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_6_0),
	.prn(vcc));
defparam \pipe[0][6] .is_wysiwyg = "true";
defparam \pipe[0][6] .power_up = "low";

dffeas \pipe[0][7] (
	.clk(clock),
	.d(\pipe~140_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~0_combout ),
	.q(pipe_7_0),
	.prn(vcc));
defparam \pipe[0][7] .is_wysiwyg = "true";
defparam \pipe[0][7] .power_up = "low";

cycloneiii_lcell_comb \pipefull~11 (
	.dataa(\pipefull[2]~q ),
	.datab(pipefull_0),
	.datac(gnd),
	.datad(accepted),
	.cin(gnd),
	.combout(\pipefull~11_combout ),
	.cout());
defparam \pipefull~11 .lut_mask = 16'hAACC;
defparam \pipefull~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_0~2 (
	.dataa(data[27]),
	.datab(data[28]),
	.datac(accepted),
	.datad(ready),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
defparam \process_0~2 .lut_mask = 16'h6996;
defparam \process_0~2 .sum_lutc_input = "datac";

dffeas \pipefull[1] (
	.clk(clock),
	.d(\pipefull~11_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~2_combout ),
	.q(\pipefull[1]~q ),
	.prn(vcc));
defparam \pipefull[1] .is_wysiwyg = "true";
defparam \pipefull[1] .power_up = "low";

cycloneiii_lcell_comb \pipefull~10 (
	.dataa(pipefull_3),
	.datab(\pipefull[1]~q ),
	.datac(gnd),
	.datad(accepted),
	.cin(gnd),
	.combout(\pipefull~10_combout ),
	.cout());
defparam \pipefull~10 .lut_mask = 16'hAACC;
defparam \pipefull~10 .sum_lutc_input = "datac";

dffeas \pipefull[2] (
	.clk(clock),
	.d(\pipefull~10_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~2_combout ),
	.q(\pipefull[2]~q ),
	.prn(vcc));
defparam \pipefull[2] .is_wysiwyg = "true";
defparam \pipefull[2] .power_up = "low";

cycloneiii_lcell_comb \pipefull[3]~9 (
	.dataa(pipefull_3),
	.datab(\pipefull[2]~q ),
	.datac(wr_en),
	.datad(gnd),
	.cin(gnd),
	.combout(\pipefull[3]~9_combout ),
	.cout());
defparam \pipefull[3]~9 .lut_mask = 16'hFEFE;
defparam \pipefull[3]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipefull[0]~12 (
	.dataa(wr_en),
	.datab(pipefull_0),
	.datac(\pipefull[1]~q ),
	.datad(accepted),
	.cin(gnd),
	.combout(\pipefull[0]~12_combout ),
	.cout());
defparam \pipefull[0]~12 .lut_mask = 16'hFEFF;
defparam \pipefull[0]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~108 (
	.dataa(\pipe[2][29]~q ),
	.datab(data[29]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~108_combout ),
	.cout());
defparam \pipe~108 .lut_mask = 16'hAACC;
defparam \pipe~108 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_1~0 (
	.dataa(accepted),
	.datab(gnd),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\process_1~0_combout ),
	.cout());
defparam \process_1~0 .lut_mask = 16'hAAFF;
defparam \process_1~0 .sum_lutc_input = "datac";

dffeas \pipe[1][29] (
	.clk(clock),
	.d(\pipe~108_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][29]~q ),
	.prn(vcc));
defparam \pipe[1][29] .is_wysiwyg = "true";
defparam \pipe[1][29] .power_up = "low";

cycloneiii_lcell_comb \pipe~90 (
	.dataa(\pipe[1][29]~q ),
	.datab(data[29]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~90_combout ),
	.cout());
defparam \pipe~90 .lut_mask = 16'hAACC;
defparam \pipe~90 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_0~0 (
	.dataa(accepted),
	.datab(gnd),
	.datac(gnd),
	.datad(pipefull_0),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
defparam \process_0~0 .lut_mask = 16'hAAFF;
defparam \process_0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~109 (
	.dataa(\pipe[2][28]~q ),
	.datab(data[28]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~109_combout ),
	.cout());
defparam \pipe~109 .lut_mask = 16'hAACC;
defparam \pipe~109 .sum_lutc_input = "datac";

dffeas \pipe[1][28] (
	.clk(clock),
	.d(\pipe~109_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][28]~q ),
	.prn(vcc));
defparam \pipe[1][28] .is_wysiwyg = "true";
defparam \pipe[1][28] .power_up = "low";

cycloneiii_lcell_comb \pipe~91 (
	.dataa(\pipe[1][28]~q ),
	.datab(data[28]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~91_combout ),
	.cout());
defparam \pipe~91 .lut_mask = 16'hAACC;
defparam \pipe~91 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~112 (
	.dataa(\pipe[2][27]~q ),
	.datab(data[27]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~112_combout ),
	.cout());
defparam \pipe~112 .lut_mask = 16'hAACC;
defparam \pipe~112 .sum_lutc_input = "datac";

dffeas \pipe[1][27] (
	.clk(clock),
	.d(\pipe~112_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][27]~q ),
	.prn(vcc));
defparam \pipe[1][27] .is_wysiwyg = "true";
defparam \pipe[1][27] .power_up = "low";

cycloneiii_lcell_comb \pipe~92 (
	.dataa(\pipe[1][27]~q ),
	.datab(data[27]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~92_combout ),
	.cout());
defparam \pipe~92 .lut_mask = 16'hAACC;
defparam \pipe~92 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~113 (
	.dataa(\pipe[2][9]~q ),
	.datab(data[9]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~113_combout ),
	.cout());
defparam \pipe~113 .lut_mask = 16'hAACC;
defparam \pipe~113 .sum_lutc_input = "datac";

dffeas \pipe[1][9] (
	.clk(clock),
	.d(\pipe~113_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][9]~q ),
	.prn(vcc));
defparam \pipe[1][9] .is_wysiwyg = "true";
defparam \pipe[1][9] .power_up = "low";

cycloneiii_lcell_comb \pipe~93 (
	.dataa(\pipe[1][9]~q ),
	.datab(data[9]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~93_combout ),
	.cout());
defparam \pipe~93 .lut_mask = 16'hAACC;
defparam \pipe~93 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~114 (
	.dataa(\pipe[2][8]~q ),
	.datab(data[8]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~114_combout ),
	.cout());
defparam \pipe~114 .lut_mask = 16'hAACC;
defparam \pipe~114 .sum_lutc_input = "datac";

dffeas \pipe[1][8] (
	.clk(clock),
	.d(\pipe~114_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][8]~q ),
	.prn(vcc));
defparam \pipe[1][8] .is_wysiwyg = "true";
defparam \pipe[1][8] .power_up = "low";

cycloneiii_lcell_comb \pipe~94 (
	.dataa(\pipe[1][8]~q ),
	.datab(data[8]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~94_combout ),
	.cout());
defparam \pipe~94 .lut_mask = 16'hAACC;
defparam \pipe~94 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~115 (
	.dataa(\pipe[2][19]~q ),
	.datab(data[19]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~115_combout ),
	.cout());
defparam \pipe~115 .lut_mask = 16'hAACC;
defparam \pipe~115 .sum_lutc_input = "datac";

dffeas \pipe[1][19] (
	.clk(clock),
	.d(\pipe~115_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][19]~q ),
	.prn(vcc));
defparam \pipe[1][19] .is_wysiwyg = "true";
defparam \pipe[1][19] .power_up = "low";

cycloneiii_lcell_comb \pipe~95 (
	.dataa(\pipe[1][19]~q ),
	.datab(data[19]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~95_combout ),
	.cout());
defparam \pipe~95 .lut_mask = 16'hAACC;
defparam \pipe~95 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~116 (
	.dataa(\pipe[2][11]~q ),
	.datab(data[11]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~116_combout ),
	.cout());
defparam \pipe~116 .lut_mask = 16'hAACC;
defparam \pipe~116 .sum_lutc_input = "datac";

dffeas \pipe[1][11] (
	.clk(clock),
	.d(\pipe~116_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][11]~q ),
	.prn(vcc));
defparam \pipe[1][11] .is_wysiwyg = "true";
defparam \pipe[1][11] .power_up = "low";

cycloneiii_lcell_comb \pipe~96 (
	.dataa(\pipe[1][11]~q ),
	.datab(data[11]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~96_combout ),
	.cout());
defparam \pipe~96 .lut_mask = 16'hAACC;
defparam \pipe~96 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~117 (
	.dataa(\pipe[2][14]~q ),
	.datab(data[14]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~117_combout ),
	.cout());
defparam \pipe~117 .lut_mask = 16'hAACC;
defparam \pipe~117 .sum_lutc_input = "datac";

dffeas \pipe[1][14] (
	.clk(clock),
	.d(\pipe~117_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][14]~q ),
	.prn(vcc));
defparam \pipe[1][14] .is_wysiwyg = "true";
defparam \pipe[1][14] .power_up = "low";

cycloneiii_lcell_comb \pipe~97 (
	.dataa(\pipe[1][14]~q ),
	.datab(data[14]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~97_combout ),
	.cout());
defparam \pipe~97 .lut_mask = 16'hAACC;
defparam \pipe~97 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~118 (
	.dataa(\pipe[2][20]~q ),
	.datab(data[20]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~118_combout ),
	.cout());
defparam \pipe~118 .lut_mask = 16'hAACC;
defparam \pipe~118 .sum_lutc_input = "datac";

dffeas \pipe[1][20] (
	.clk(clock),
	.d(\pipe~118_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][20]~q ),
	.prn(vcc));
defparam \pipe[1][20] .is_wysiwyg = "true";
defparam \pipe[1][20] .power_up = "low";

cycloneiii_lcell_comb \pipe~98 (
	.dataa(\pipe[1][20]~q ),
	.datab(data[20]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~98_combout ),
	.cout());
defparam \pipe~98 .lut_mask = 16'hAACC;
defparam \pipe~98 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~119 (
	.dataa(\pipe[2][18]~q ),
	.datab(data[18]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~119_combout ),
	.cout());
defparam \pipe~119 .lut_mask = 16'hAACC;
defparam \pipe~119 .sum_lutc_input = "datac";

dffeas \pipe[1][18] (
	.clk(clock),
	.d(\pipe~119_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][18]~q ),
	.prn(vcc));
defparam \pipe[1][18] .is_wysiwyg = "true";
defparam \pipe[1][18] .power_up = "low";

cycloneiii_lcell_comb \pipe~99 (
	.dataa(\pipe[1][18]~q ),
	.datab(data[18]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~99_combout ),
	.cout());
defparam \pipe~99 .lut_mask = 16'hAACC;
defparam \pipe~99 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~120 (
	.dataa(\pipe[2][13]~q ),
	.datab(data[13]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~120_combout ),
	.cout());
defparam \pipe~120 .lut_mask = 16'hAACC;
defparam \pipe~120 .sum_lutc_input = "datac";

dffeas \pipe[1][13] (
	.clk(clock),
	.d(\pipe~120_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][13]~q ),
	.prn(vcc));
defparam \pipe[1][13] .is_wysiwyg = "true";
defparam \pipe[1][13] .power_up = "low";

cycloneiii_lcell_comb \pipe~100 (
	.dataa(\pipe[1][13]~q ),
	.datab(data[13]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~100_combout ),
	.cout());
defparam \pipe~100 .lut_mask = 16'hAACC;
defparam \pipe~100 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~121 (
	.dataa(\pipe[2][15]~q ),
	.datab(data[15]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~121_combout ),
	.cout());
defparam \pipe~121 .lut_mask = 16'hAACC;
defparam \pipe~121 .sum_lutc_input = "datac";

dffeas \pipe[1][15] (
	.clk(clock),
	.d(\pipe~121_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][15]~q ),
	.prn(vcc));
defparam \pipe[1][15] .is_wysiwyg = "true";
defparam \pipe[1][15] .power_up = "low";

cycloneiii_lcell_comb \pipe~101 (
	.dataa(\pipe[1][15]~q ),
	.datab(data[15]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~101_combout ),
	.cout());
defparam \pipe~101 .lut_mask = 16'hAACC;
defparam \pipe~101 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~122 (
	.dataa(\pipe[2][10]~q ),
	.datab(data[10]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~122_combout ),
	.cout());
defparam \pipe~122 .lut_mask = 16'hAACC;
defparam \pipe~122 .sum_lutc_input = "datac";

dffeas \pipe[1][10] (
	.clk(clock),
	.d(\pipe~122_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][10]~q ),
	.prn(vcc));
defparam \pipe[1][10] .is_wysiwyg = "true";
defparam \pipe[1][10] .power_up = "low";

cycloneiii_lcell_comb \pipe~102 (
	.dataa(\pipe[1][10]~q ),
	.datab(data[10]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~102_combout ),
	.cout());
defparam \pipe~102 .lut_mask = 16'hAACC;
defparam \pipe~102 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~123 (
	.dataa(\pipe[2][16]~q ),
	.datab(data[16]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~123_combout ),
	.cout());
defparam \pipe~123 .lut_mask = 16'hAACC;
defparam \pipe~123 .sum_lutc_input = "datac";

dffeas \pipe[1][16] (
	.clk(clock),
	.d(\pipe~123_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][16]~q ),
	.prn(vcc));
defparam \pipe[1][16] .is_wysiwyg = "true";
defparam \pipe[1][16] .power_up = "low";

cycloneiii_lcell_comb \pipe~103 (
	.dataa(\pipe[1][16]~q ),
	.datab(data[16]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~103_combout ),
	.cout());
defparam \pipe~103 .lut_mask = 16'hAACC;
defparam \pipe~103 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~124 (
	.dataa(\pipe[2][17]~q ),
	.datab(data[17]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~124_combout ),
	.cout());
defparam \pipe~124 .lut_mask = 16'hAACC;
defparam \pipe~124 .sum_lutc_input = "datac";

dffeas \pipe[1][17] (
	.clk(clock),
	.d(\pipe~124_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][17]~q ),
	.prn(vcc));
defparam \pipe[1][17] .is_wysiwyg = "true";
defparam \pipe[1][17] .power_up = "low";

cycloneiii_lcell_comb \pipe~104 (
	.dataa(\pipe[1][17]~q ),
	.datab(data[17]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~104_combout ),
	.cout());
defparam \pipe~104 .lut_mask = 16'hAACC;
defparam \pipe~104 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~125 (
	.dataa(\pipe[2][21]~q ),
	.datab(data[21]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~125_combout ),
	.cout());
defparam \pipe~125 .lut_mask = 16'hAACC;
defparam \pipe~125 .sum_lutc_input = "datac";

dffeas \pipe[1][21] (
	.clk(clock),
	.d(\pipe~125_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][21]~q ),
	.prn(vcc));
defparam \pipe[1][21] .is_wysiwyg = "true";
defparam \pipe[1][21] .power_up = "low";

cycloneiii_lcell_comb \pipe~105 (
	.dataa(\pipe[1][21]~q ),
	.datab(data[21]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~105_combout ),
	.cout());
defparam \pipe~105 .lut_mask = 16'hAACC;
defparam \pipe~105 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~126 (
	.dataa(\pipe[2][12]~q ),
	.datab(data[12]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~126_combout ),
	.cout());
defparam \pipe~126 .lut_mask = 16'hAACC;
defparam \pipe~126 .sum_lutc_input = "datac";

dffeas \pipe[1][12] (
	.clk(clock),
	.d(\pipe~126_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][12]~q ),
	.prn(vcc));
defparam \pipe[1][12] .is_wysiwyg = "true";
defparam \pipe[1][12] .power_up = "low";

cycloneiii_lcell_comb \pipe~106 (
	.dataa(\pipe[1][12]~q ),
	.datab(data[12]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~106_combout ),
	.cout());
defparam \pipe~106 .lut_mask = 16'hAACC;
defparam \pipe~106 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~127 (
	.dataa(\pipe[2][22]~q ),
	.datab(data[22]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~127_combout ),
	.cout());
defparam \pipe~127 .lut_mask = 16'hAACC;
defparam \pipe~127 .sum_lutc_input = "datac";

dffeas \pipe[1][22] (
	.clk(clock),
	.d(\pipe~127_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][22]~q ),
	.prn(vcc));
defparam \pipe[1][22] .is_wysiwyg = "true";
defparam \pipe[1][22] .power_up = "low";

cycloneiii_lcell_comb \pipe~107 (
	.dataa(\pipe[1][22]~q ),
	.datab(data[22]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~107_combout ),
	.cout());
defparam \pipe~107 .lut_mask = 16'hAACC;
defparam \pipe~107 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~130 (
	.dataa(\pipe[2][24]~q ),
	.datab(data[24]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~130_combout ),
	.cout());
defparam \pipe~130 .lut_mask = 16'hAACC;
defparam \pipe~130 .sum_lutc_input = "datac";

dffeas \pipe[1][24] (
	.clk(clock),
	.d(\pipe~130_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][24]~q ),
	.prn(vcc));
defparam \pipe[1][24] .is_wysiwyg = "true";
defparam \pipe[1][24] .power_up = "low";

cycloneiii_lcell_comb \pipe~110 (
	.dataa(\pipe[1][24]~q ),
	.datab(data[24]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~110_combout ),
	.cout());
defparam \pipe~110 .lut_mask = 16'hAACC;
defparam \pipe~110 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~131 (
	.dataa(\pipe[2][25]~q ),
	.datab(data[25]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~131_combout ),
	.cout());
defparam \pipe~131 .lut_mask = 16'hAACC;
defparam \pipe~131 .sum_lutc_input = "datac";

dffeas \pipe[1][25] (
	.clk(clock),
	.d(\pipe~131_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][25]~q ),
	.prn(vcc));
defparam \pipe[1][25] .is_wysiwyg = "true";
defparam \pipe[1][25] .power_up = "low";

cycloneiii_lcell_comb \pipe~111 (
	.dataa(\pipe[1][25]~q ),
	.datab(data[25]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~111_combout ),
	.cout());
defparam \pipe~111 .lut_mask = 16'hAACC;
defparam \pipe~111 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~158 (
	.dataa(\pipe[2][0]~q ),
	.datab(data[0]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~158_combout ),
	.cout());
defparam \pipe~158 .lut_mask = 16'hAACC;
defparam \pipe~158 .sum_lutc_input = "datac";

dffeas \pipe[1][0] (
	.clk(clock),
	.d(\pipe~158_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][0]~q ),
	.prn(vcc));
defparam \pipe[1][0] .is_wysiwyg = "true";
defparam \pipe[1][0] .power_up = "low";

cycloneiii_lcell_comb \pipe~133 (
	.dataa(\pipe[1][0]~q ),
	.datab(data[0]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~133_combout ),
	.cout());
defparam \pipe~133 .lut_mask = 16'hAACC;
defparam \pipe~133 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~159 (
	.dataa(\pipe[2][1]~q ),
	.datab(data[1]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~159_combout ),
	.cout());
defparam \pipe~159 .lut_mask = 16'hAACC;
defparam \pipe~159 .sum_lutc_input = "datac";

dffeas \pipe[1][1] (
	.clk(clock),
	.d(\pipe~159_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][1]~q ),
	.prn(vcc));
defparam \pipe[1][1] .is_wysiwyg = "true";
defparam \pipe[1][1] .power_up = "low";

cycloneiii_lcell_comb \pipe~134 (
	.dataa(\pipe[1][1]~q ),
	.datab(data[1]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~134_combout ),
	.cout());
defparam \pipe~134 .lut_mask = 16'hAACC;
defparam \pipe~134 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~160 (
	.dataa(\pipe[2][2]~q ),
	.datab(data[2]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~160_combout ),
	.cout());
defparam \pipe~160 .lut_mask = 16'hAACC;
defparam \pipe~160 .sum_lutc_input = "datac";

dffeas \pipe[1][2] (
	.clk(clock),
	.d(\pipe~160_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][2]~q ),
	.prn(vcc));
defparam \pipe[1][2] .is_wysiwyg = "true";
defparam \pipe[1][2] .power_up = "low";

cycloneiii_lcell_comb \pipe~135 (
	.dataa(\pipe[1][2]~q ),
	.datab(data[2]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~135_combout ),
	.cout());
defparam \pipe~135 .lut_mask = 16'hAACC;
defparam \pipe~135 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~161 (
	.dataa(\pipe[2][3]~q ),
	.datab(data[3]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~161_combout ),
	.cout());
defparam \pipe~161 .lut_mask = 16'hAACC;
defparam \pipe~161 .sum_lutc_input = "datac";

dffeas \pipe[1][3] (
	.clk(clock),
	.d(\pipe~161_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][3]~q ),
	.prn(vcc));
defparam \pipe[1][3] .is_wysiwyg = "true";
defparam \pipe[1][3] .power_up = "low";

cycloneiii_lcell_comb \pipe~136 (
	.dataa(\pipe[1][3]~q ),
	.datab(data[3]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~136_combout ),
	.cout());
defparam \pipe~136 .lut_mask = 16'hAACC;
defparam \pipe~136 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~162 (
	.dataa(\pipe[2][4]~q ),
	.datab(data[4]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~162_combout ),
	.cout());
defparam \pipe~162 .lut_mask = 16'hAACC;
defparam \pipe~162 .sum_lutc_input = "datac";

dffeas \pipe[1][4] (
	.clk(clock),
	.d(\pipe~162_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][4]~q ),
	.prn(vcc));
defparam \pipe[1][4] .is_wysiwyg = "true";
defparam \pipe[1][4] .power_up = "low";

cycloneiii_lcell_comb \pipe~137 (
	.dataa(\pipe[1][4]~q ),
	.datab(data[4]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~137_combout ),
	.cout());
defparam \pipe~137 .lut_mask = 16'hAACC;
defparam \pipe~137 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~163 (
	.dataa(\pipe[2][5]~q ),
	.datab(data[5]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~163_combout ),
	.cout());
defparam \pipe~163 .lut_mask = 16'hAACC;
defparam \pipe~163 .sum_lutc_input = "datac";

dffeas \pipe[1][5] (
	.clk(clock),
	.d(\pipe~163_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][5]~q ),
	.prn(vcc));
defparam \pipe[1][5] .is_wysiwyg = "true";
defparam \pipe[1][5] .power_up = "low";

cycloneiii_lcell_comb \pipe~138 (
	.dataa(\pipe[1][5]~q ),
	.datab(data[5]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~138_combout ),
	.cout());
defparam \pipe~138 .lut_mask = 16'hAACC;
defparam \pipe~138 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~164 (
	.dataa(\pipe[2][6]~q ),
	.datab(data[6]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~164_combout ),
	.cout());
defparam \pipe~164 .lut_mask = 16'hAACC;
defparam \pipe~164 .sum_lutc_input = "datac";

dffeas \pipe[1][6] (
	.clk(clock),
	.d(\pipe~164_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][6]~q ),
	.prn(vcc));
defparam \pipe[1][6] .is_wysiwyg = "true";
defparam \pipe[1][6] .power_up = "low";

cycloneiii_lcell_comb \pipe~139 (
	.dataa(\pipe[1][6]~q ),
	.datab(data[6]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~139_combout ),
	.cout());
defparam \pipe~139 .lut_mask = 16'hAACC;
defparam \pipe~139 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pipe~165 (
	.dataa(\pipe[2][7]~q ),
	.datab(data[7]),
	.datac(gnd),
	.datad(\pipefull[2]~q ),
	.cin(gnd),
	.combout(\pipe~165_combout ),
	.cout());
defparam \pipe~165 .lut_mask = 16'hAACC;
defparam \pipe~165 .sum_lutc_input = "datac";

dffeas \pipe[1][7] (
	.clk(clock),
	.d(\pipe~165_combout ),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_1~0_combout ),
	.q(\pipe[1][7]~q ),
	.prn(vcc));
defparam \pipe[1][7] .is_wysiwyg = "true";
defparam \pipe[1][7] .power_up = "low";

cycloneiii_lcell_comb \pipe~140 (
	.dataa(\pipe[1][7]~q ),
	.datab(data[7]),
	.datac(gnd),
	.datad(\pipefull[1]~q ),
	.cin(gnd),
	.combout(\pipe~140_combout ),
	.cout());
defparam \pipe~140 .lut_mask = 16'hAACC;
defparam \pipe~140 .sum_lutc_input = "datac";

endmodule

module altera_ddr_auk_ddr_hp_timers (
	clk,
	reset_n,
	am_writing,
	doing_act,
	twr_pipe_2,
	to_this_bank_0,
	finished_twr1,
	finished_tras1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	am_writing;
input 	doing_act;
output 	twr_pipe_2;
input 	to_this_bank_0;
output 	finished_twr1;
output 	finished_tras1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \tras_pipe[1]~q ;
wire \tras_pipe[0]~q ;
wire \tras_pipe~16_combout ;
wire \start_ap_trcd_timer~combout ;
wire \start_twr_timer~combout ;
wire \twr_pipe[0]~q ;
wire \twr_pipe~7_combout ;
wire \twr_pipe[1]~q ;
wire \twr_pipe~6_combout ;
wire \tras_pipe~15_combout ;
wire \tras_pipe[2]~q ;


dffeas \tras_pipe[1] (
	.clk(clk),
	.d(\tras_pipe~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[1]~q ),
	.prn(vcc));
defparam \tras_pipe[1] .is_wysiwyg = "true";
defparam \tras_pipe[1] .power_up = "low";

dffeas \tras_pipe[0] (
	.clk(clk),
	.d(\start_ap_trcd_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[0]~q ),
	.prn(vcc));
defparam \tras_pipe[0] .is_wysiwyg = "true";
defparam \tras_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \tras_pipe~16 (
	.dataa(\tras_pipe[0]~q ),
	.datab(to_this_bank_0),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~16_combout ),
	.cout());
defparam \tras_pipe~16 .lut_mask = 16'hEEFF;
defparam \tras_pipe~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb start_ap_trcd_timer(
	.dataa(doing_act),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_0),
	.cin(gnd),
	.combout(\start_ap_trcd_timer~combout ),
	.cout());
defparam start_ap_trcd_timer.lut_mask = 16'hFF55;
defparam start_ap_trcd_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[2] (
	.clk(clk),
	.d(\twr_pipe~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(twr_pipe_2),
	.prn(vcc));
defparam \twr_pipe[2] .is_wysiwyg = "true";
defparam \twr_pipe[2] .power_up = "low";

cycloneiii_lcell_comb finished_twr(
	.dataa(to_this_bank_0),
	.datab(gnd),
	.datac(am_writing),
	.datad(twr_pipe_2),
	.cin(gnd),
	.combout(finished_twr1),
	.cout());
defparam finished_twr.lut_mask = 16'hAFFF;
defparam finished_twr.sum_lutc_input = "datac";

dffeas finished_tras(
	.clk(clk),
	.d(\tras_pipe[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(finished_tras1),
	.prn(vcc));
defparam finished_tras.is_wysiwyg = "true";
defparam finished_tras.power_up = "low";

cycloneiii_lcell_comb start_twr_timer(
	.dataa(am_writing),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_0),
	.cin(gnd),
	.combout(\start_twr_timer~combout ),
	.cout());
defparam start_twr_timer.lut_mask = 16'hAAFF;
defparam start_twr_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[0] (
	.clk(clk),
	.d(\start_twr_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[0]~q ),
	.prn(vcc));
defparam \twr_pipe[0] .is_wysiwyg = "true";
defparam \twr_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~7 (
	.dataa(to_this_bank_0),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[0]~q ),
	.cin(gnd),
	.combout(\twr_pipe~7_combout ),
	.cout());
defparam \twr_pipe~7 .lut_mask = 16'hFFF5;
defparam \twr_pipe~7 .sum_lutc_input = "datac";

dffeas \twr_pipe[1] (
	.clk(clk),
	.d(\twr_pipe~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[1]~q ),
	.prn(vcc));
defparam \twr_pipe[1] .is_wysiwyg = "true";
defparam \twr_pipe[1] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~6 (
	.dataa(to_this_bank_0),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[1]~q ),
	.cin(gnd),
	.combout(\twr_pipe~6_combout ),
	.cout());
defparam \twr_pipe~6 .lut_mask = 16'hFFF5;
defparam \twr_pipe~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tras_pipe~15 (
	.dataa(\tras_pipe[1]~q ),
	.datab(to_this_bank_0),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~15_combout ),
	.cout());
defparam \tras_pipe~15 .lut_mask = 16'hEEFF;
defparam \tras_pipe~15 .sum_lutc_input = "datac";

dffeas \tras_pipe[2] (
	.clk(clk),
	.d(\tras_pipe~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[2]~q ),
	.prn(vcc));
defparam \tras_pipe[2] .is_wysiwyg = "true";
defparam \tras_pipe[2] .power_up = "low";

endmodule

module altera_ddr_auk_ddr_hp_timers_1 (
	clk,
	reset_n,
	am_writing,
	doing_act,
	twr_pipe_2,
	to_this_bank_1,
	finished_twr1,
	finished_tras1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	am_writing;
input 	doing_act;
output 	twr_pipe_2;
input 	to_this_bank_1;
output 	finished_twr1;
output 	finished_tras1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \tras_pipe[1]~q ;
wire \tras_pipe[0]~q ;
wire \tras_pipe~16_combout ;
wire \start_ap_trcd_timer~combout ;
wire \start_twr_timer~combout ;
wire \twr_pipe[0]~q ;
wire \twr_pipe~7_combout ;
wire \twr_pipe[1]~q ;
wire \twr_pipe~6_combout ;
wire \tras_pipe~15_combout ;
wire \tras_pipe[2]~q ;


dffeas \tras_pipe[1] (
	.clk(clk),
	.d(\tras_pipe~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[1]~q ),
	.prn(vcc));
defparam \tras_pipe[1] .is_wysiwyg = "true";
defparam \tras_pipe[1] .power_up = "low";

dffeas \tras_pipe[0] (
	.clk(clk),
	.d(\start_ap_trcd_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[0]~q ),
	.prn(vcc));
defparam \tras_pipe[0] .is_wysiwyg = "true";
defparam \tras_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \tras_pipe~16 (
	.dataa(\tras_pipe[0]~q ),
	.datab(to_this_bank_1),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~16_combout ),
	.cout());
defparam \tras_pipe~16 .lut_mask = 16'hEEFF;
defparam \tras_pipe~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb start_ap_trcd_timer(
	.dataa(doing_act),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_1),
	.cin(gnd),
	.combout(\start_ap_trcd_timer~combout ),
	.cout());
defparam start_ap_trcd_timer.lut_mask = 16'hFF55;
defparam start_ap_trcd_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[2] (
	.clk(clk),
	.d(\twr_pipe~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(twr_pipe_2),
	.prn(vcc));
defparam \twr_pipe[2] .is_wysiwyg = "true";
defparam \twr_pipe[2] .power_up = "low";

cycloneiii_lcell_comb finished_twr(
	.dataa(to_this_bank_1),
	.datab(gnd),
	.datac(am_writing),
	.datad(twr_pipe_2),
	.cin(gnd),
	.combout(finished_twr1),
	.cout());
defparam finished_twr.lut_mask = 16'hAFFF;
defparam finished_twr.sum_lutc_input = "datac";

dffeas finished_tras(
	.clk(clk),
	.d(\tras_pipe[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(finished_tras1),
	.prn(vcc));
defparam finished_tras.is_wysiwyg = "true";
defparam finished_tras.power_up = "low";

cycloneiii_lcell_comb start_twr_timer(
	.dataa(am_writing),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_1),
	.cin(gnd),
	.combout(\start_twr_timer~combout ),
	.cout());
defparam start_twr_timer.lut_mask = 16'hAAFF;
defparam start_twr_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[0] (
	.clk(clk),
	.d(\start_twr_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[0]~q ),
	.prn(vcc));
defparam \twr_pipe[0] .is_wysiwyg = "true";
defparam \twr_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~7 (
	.dataa(to_this_bank_1),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[0]~q ),
	.cin(gnd),
	.combout(\twr_pipe~7_combout ),
	.cout());
defparam \twr_pipe~7 .lut_mask = 16'hFFF5;
defparam \twr_pipe~7 .sum_lutc_input = "datac";

dffeas \twr_pipe[1] (
	.clk(clk),
	.d(\twr_pipe~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[1]~q ),
	.prn(vcc));
defparam \twr_pipe[1] .is_wysiwyg = "true";
defparam \twr_pipe[1] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~6 (
	.dataa(to_this_bank_1),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[1]~q ),
	.cin(gnd),
	.combout(\twr_pipe~6_combout ),
	.cout());
defparam \twr_pipe~6 .lut_mask = 16'hFFF5;
defparam \twr_pipe~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tras_pipe~15 (
	.dataa(\tras_pipe[1]~q ),
	.datab(to_this_bank_1),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~15_combout ),
	.cout());
defparam \tras_pipe~15 .lut_mask = 16'hEEFF;
defparam \tras_pipe~15 .sum_lutc_input = "datac";

dffeas \tras_pipe[2] (
	.clk(clk),
	.d(\tras_pipe~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[2]~q ),
	.prn(vcc));
defparam \tras_pipe[2] .is_wysiwyg = "true";
defparam \tras_pipe[2] .power_up = "low";

endmodule

module altera_ddr_auk_ddr_hp_timers_2 (
	clk,
	reset_n,
	am_writing,
	doing_act,
	twr_pipe_2,
	to_this_bank_2,
	finished_twr1,
	finished_tras1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	am_writing;
input 	doing_act;
output 	twr_pipe_2;
input 	to_this_bank_2;
output 	finished_twr1;
output 	finished_tras1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \tras_pipe[1]~q ;
wire \tras_pipe[0]~q ;
wire \tras_pipe~16_combout ;
wire \start_ap_trcd_timer~combout ;
wire \start_twr_timer~combout ;
wire \twr_pipe[0]~q ;
wire \twr_pipe~7_combout ;
wire \twr_pipe[1]~q ;
wire \twr_pipe~6_combout ;
wire \tras_pipe~15_combout ;
wire \tras_pipe[2]~q ;


dffeas \tras_pipe[1] (
	.clk(clk),
	.d(\tras_pipe~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[1]~q ),
	.prn(vcc));
defparam \tras_pipe[1] .is_wysiwyg = "true";
defparam \tras_pipe[1] .power_up = "low";

dffeas \tras_pipe[0] (
	.clk(clk),
	.d(\start_ap_trcd_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[0]~q ),
	.prn(vcc));
defparam \tras_pipe[0] .is_wysiwyg = "true";
defparam \tras_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \tras_pipe~16 (
	.dataa(\tras_pipe[0]~q ),
	.datab(to_this_bank_2),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~16_combout ),
	.cout());
defparam \tras_pipe~16 .lut_mask = 16'hEEFF;
defparam \tras_pipe~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb start_ap_trcd_timer(
	.dataa(doing_act),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_2),
	.cin(gnd),
	.combout(\start_ap_trcd_timer~combout ),
	.cout());
defparam start_ap_trcd_timer.lut_mask = 16'hFF55;
defparam start_ap_trcd_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[2] (
	.clk(clk),
	.d(\twr_pipe~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(twr_pipe_2),
	.prn(vcc));
defparam \twr_pipe[2] .is_wysiwyg = "true";
defparam \twr_pipe[2] .power_up = "low";

cycloneiii_lcell_comb finished_twr(
	.dataa(to_this_bank_2),
	.datab(gnd),
	.datac(am_writing),
	.datad(twr_pipe_2),
	.cin(gnd),
	.combout(finished_twr1),
	.cout());
defparam finished_twr.lut_mask = 16'hAFFF;
defparam finished_twr.sum_lutc_input = "datac";

dffeas finished_tras(
	.clk(clk),
	.d(\tras_pipe[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(finished_tras1),
	.prn(vcc));
defparam finished_tras.is_wysiwyg = "true";
defparam finished_tras.power_up = "low";

cycloneiii_lcell_comb start_twr_timer(
	.dataa(am_writing),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_2),
	.cin(gnd),
	.combout(\start_twr_timer~combout ),
	.cout());
defparam start_twr_timer.lut_mask = 16'hAAFF;
defparam start_twr_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[0] (
	.clk(clk),
	.d(\start_twr_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[0]~q ),
	.prn(vcc));
defparam \twr_pipe[0] .is_wysiwyg = "true";
defparam \twr_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~7 (
	.dataa(to_this_bank_2),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[0]~q ),
	.cin(gnd),
	.combout(\twr_pipe~7_combout ),
	.cout());
defparam \twr_pipe~7 .lut_mask = 16'hFFF5;
defparam \twr_pipe~7 .sum_lutc_input = "datac";

dffeas \twr_pipe[1] (
	.clk(clk),
	.d(\twr_pipe~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[1]~q ),
	.prn(vcc));
defparam \twr_pipe[1] .is_wysiwyg = "true";
defparam \twr_pipe[1] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~6 (
	.dataa(to_this_bank_2),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[1]~q ),
	.cin(gnd),
	.combout(\twr_pipe~6_combout ),
	.cout());
defparam \twr_pipe~6 .lut_mask = 16'hFFF5;
defparam \twr_pipe~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tras_pipe~15 (
	.dataa(\tras_pipe[1]~q ),
	.datab(to_this_bank_2),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~15_combout ),
	.cout());
defparam \tras_pipe~15 .lut_mask = 16'hEEFF;
defparam \tras_pipe~15 .sum_lutc_input = "datac";

dffeas \tras_pipe[2] (
	.clk(clk),
	.d(\tras_pipe~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[2]~q ),
	.prn(vcc));
defparam \tras_pipe[2] .is_wysiwyg = "true";
defparam \tras_pipe[2] .power_up = "low";

endmodule

module altera_ddr_auk_ddr_hp_timers_3 (
	clk,
	reset_n,
	am_writing,
	doing_act,
	twr_pipe_2,
	to_this_bank_3,
	finished_twr1,
	finished_tras1)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	reset_n;
input 	am_writing;
input 	doing_act;
output 	twr_pipe_2;
input 	to_this_bank_3;
output 	finished_twr1;
output 	finished_tras1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \tras_pipe[1]~q ;
wire \tras_pipe[0]~q ;
wire \tras_pipe~16_combout ;
wire \start_ap_trcd_timer~combout ;
wire \start_twr_timer~combout ;
wire \twr_pipe[0]~q ;
wire \twr_pipe~7_combout ;
wire \twr_pipe[1]~q ;
wire \twr_pipe~6_combout ;
wire \tras_pipe~15_combout ;
wire \tras_pipe[2]~q ;


dffeas \tras_pipe[1] (
	.clk(clk),
	.d(\tras_pipe~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[1]~q ),
	.prn(vcc));
defparam \tras_pipe[1] .is_wysiwyg = "true";
defparam \tras_pipe[1] .power_up = "low";

dffeas \tras_pipe[0] (
	.clk(clk),
	.d(\start_ap_trcd_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[0]~q ),
	.prn(vcc));
defparam \tras_pipe[0] .is_wysiwyg = "true";
defparam \tras_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \tras_pipe~16 (
	.dataa(\tras_pipe[0]~q ),
	.datab(to_this_bank_3),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~16_combout ),
	.cout());
defparam \tras_pipe~16 .lut_mask = 16'hEEFF;
defparam \tras_pipe~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb start_ap_trcd_timer(
	.dataa(doing_act),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_3),
	.cin(gnd),
	.combout(\start_ap_trcd_timer~combout ),
	.cout());
defparam start_ap_trcd_timer.lut_mask = 16'hFF55;
defparam start_ap_trcd_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[2] (
	.clk(clk),
	.d(\twr_pipe~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(twr_pipe_2),
	.prn(vcc));
defparam \twr_pipe[2] .is_wysiwyg = "true";
defparam \twr_pipe[2] .power_up = "low";

cycloneiii_lcell_comb finished_twr(
	.dataa(to_this_bank_3),
	.datab(gnd),
	.datac(am_writing),
	.datad(twr_pipe_2),
	.cin(gnd),
	.combout(finished_twr1),
	.cout());
defparam finished_twr.lut_mask = 16'hAFFF;
defparam finished_twr.sum_lutc_input = "datac";

dffeas finished_tras(
	.clk(clk),
	.d(\tras_pipe[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(finished_tras1),
	.prn(vcc));
defparam finished_tras.is_wysiwyg = "true";
defparam finished_tras.power_up = "low";

cycloneiii_lcell_comb start_twr_timer(
	.dataa(am_writing),
	.datab(gnd),
	.datac(gnd),
	.datad(to_this_bank_3),
	.cin(gnd),
	.combout(\start_twr_timer~combout ),
	.cout());
defparam start_twr_timer.lut_mask = 16'hAAFF;
defparam start_twr_timer.sum_lutc_input = "datac";

dffeas \twr_pipe[0] (
	.clk(clk),
	.d(\start_twr_timer~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[0]~q ),
	.prn(vcc));
defparam \twr_pipe[0] .is_wysiwyg = "true";
defparam \twr_pipe[0] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~7 (
	.dataa(to_this_bank_3),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[0]~q ),
	.cin(gnd),
	.combout(\twr_pipe~7_combout ),
	.cout());
defparam \twr_pipe~7 .lut_mask = 16'hFFF5;
defparam \twr_pipe~7 .sum_lutc_input = "datac";

dffeas \twr_pipe[1] (
	.clk(clk),
	.d(\twr_pipe~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\twr_pipe[1]~q ),
	.prn(vcc));
defparam \twr_pipe[1] .is_wysiwyg = "true";
defparam \twr_pipe[1] .power_up = "low";

cycloneiii_lcell_comb \twr_pipe~6 (
	.dataa(to_this_bank_3),
	.datab(gnd),
	.datac(am_writing),
	.datad(\twr_pipe[1]~q ),
	.cin(gnd),
	.combout(\twr_pipe~6_combout ),
	.cout());
defparam \twr_pipe~6 .lut_mask = 16'hFFF5;
defparam \twr_pipe~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tras_pipe~15 (
	.dataa(\tras_pipe[1]~q ),
	.datab(to_this_bank_3),
	.datac(gnd),
	.datad(doing_act),
	.cin(gnd),
	.combout(\tras_pipe~15_combout ),
	.cout());
defparam \tras_pipe~15 .lut_mask = 16'hEEFF;
defparam \tras_pipe~15 .sum_lutc_input = "datac";

dffeas \tras_pipe[2] (
	.clk(clk),
	.d(\tras_pipe~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tras_pipe[2]~q ),
	.prn(vcc));
defparam \tras_pipe[2] .is_wysiwyg = "true";
defparam \tras_pipe[2] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy (
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dm_ddio_dataout_0,
	dm_ddio_dataout_1,
	ddio_outa_0,
	ddio_outa_01,
	dq_ddio_dataout_0,
	dq_ddio_dataout_1,
	dq_ddio_dataout_2,
	dq_ddio_dataout_3,
	dq_ddio_dataout_4,
	dq_ddio_dataout_5,
	dq_ddio_dataout_6,
	dq_ddio_dataout_7,
	dq_ddio_dataout_8,
	dq_ddio_dataout_9,
	dq_ddio_dataout_10,
	dq_ddio_dataout_11,
	dq_ddio_dataout_12,
	dq_ddio_dataout_13,
	dq_ddio_dataout_14,
	dq_ddio_dataout_15,
	dqs_ddio_dataout_0,
	wdp_wdqs_oe_2x_r_0,
	dqs_ddio_dataout_1,
	wdp_wdqs_oe_2x_r_1,
	q_b_34,
	q_b_32,
	q_b_35,
	q_b_33,
	q_b_161,
	q_b_01,
	q_b_171,
	q_b_110,
	q_b_181,
	q_b_210,
	q_b_191,
	q_b_36,
	q_b_201,
	q_b_41,
	q_b_211,
	q_b_51,
	q_b_221,
	q_b_61,
	q_b_231,
	q_b_71,
	q_b_241,
	q_b_81,
	q_b_251,
	q_b_91,
	q_b_261,
	q_b_101,
	q_b_271,
	q_b_111,
	q_b_281,
	q_b_121,
	q_b_291,
	q_b_131,
	q_b_301,
	q_b_141,
	q_b_311,
	q_b_151,
	seq_ac_add_1t_ac_lat_internal,
	ctl_rdata_valid_0,
	reset_request_n,
	ctl_init_success,
	reset_phy_clk_1x_n,
	control_doing_rd_0,
	cs_n_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	ba_0,
	ba_1,
	ras_n,
	cas_n,
	we_n,
	wdp_wdata_oe_2x_r_0,
	wdp_wdata_oe_2x_r_1,
	wdp_wdata_oe_2x_r_2,
	wdp_wdata_oe_2x_r_3,
	wdp_wdata_oe_2x_r_4,
	wdp_wdata_oe_2x_r_5,
	wdp_wdata_oe_2x_r_6,
	wdp_wdata_oe_2x_r_7,
	wdp_wdata_oe_2x_r_8,
	wdp_wdata_oe_2x_r_9,
	wdp_wdata_oe_2x_r_10,
	wdp_wdata_oe_2x_r_11,
	wdp_wdata_oe_2x_r_12,
	wdp_wdata_oe_2x_r_13,
	wdp_wdata_oe_2x_r_14,
	wdp_wdata_oe_2x_r_15,
	control_wlat_r_0,
	control_doing_wr,
	Equal6,
	control_doing_wr1,
	control_doing_wr2,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	control_dqs_burst_0,
	dqs_burst_cas4,
	dqs_burst_cas3,
	GND_port,
	mem_clk_0,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=1 */;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dm_ddio_dataout_0;
output 	dm_ddio_dataout_1;
output 	ddio_outa_0;
output 	ddio_outa_01;
output 	dq_ddio_dataout_0;
output 	dq_ddio_dataout_1;
output 	dq_ddio_dataout_2;
output 	dq_ddio_dataout_3;
output 	dq_ddio_dataout_4;
output 	dq_ddio_dataout_5;
output 	dq_ddio_dataout_6;
output 	dq_ddio_dataout_7;
output 	dq_ddio_dataout_8;
output 	dq_ddio_dataout_9;
output 	dq_ddio_dataout_10;
output 	dq_ddio_dataout_11;
output 	dq_ddio_dataout_12;
output 	dq_ddio_dataout_13;
output 	dq_ddio_dataout_14;
output 	dq_ddio_dataout_15;
output 	dqs_ddio_dataout_0;
output 	wdp_wdqs_oe_2x_r_0;
output 	dqs_ddio_dataout_1;
output 	wdp_wdqs_oe_2x_r_1;
input 	q_b_34;
input 	q_b_32;
input 	q_b_35;
input 	q_b_33;
input 	q_b_161;
input 	q_b_01;
input 	q_b_171;
input 	q_b_110;
input 	q_b_181;
input 	q_b_210;
input 	q_b_191;
input 	q_b_36;
input 	q_b_201;
input 	q_b_41;
input 	q_b_211;
input 	q_b_51;
input 	q_b_221;
input 	q_b_61;
input 	q_b_231;
input 	q_b_71;
input 	q_b_241;
input 	q_b_81;
input 	q_b_251;
input 	q_b_91;
input 	q_b_261;
input 	q_b_101;
input 	q_b_271;
input 	q_b_111;
input 	q_b_281;
input 	q_b_121;
input 	q_b_291;
input 	q_b_131;
input 	q_b_301;
input 	q_b_141;
input 	q_b_311;
input 	q_b_151;
output 	seq_ac_add_1t_ac_lat_internal;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	ctl_init_success;
output 	reset_phy_clk_1x_n;
input 	control_doing_rd_0;
input 	cs_n_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	ba_0;
input 	ba_1;
input 	ras_n;
input 	cas_n;
input 	we_n;
output 	wdp_wdata_oe_2x_r_0;
output 	wdp_wdata_oe_2x_r_1;
output 	wdp_wdata_oe_2x_r_2;
output 	wdp_wdata_oe_2x_r_3;
output 	wdp_wdata_oe_2x_r_4;
output 	wdp_wdata_oe_2x_r_5;
output 	wdp_wdata_oe_2x_r_6;
output 	wdp_wdata_oe_2x_r_7;
output 	wdp_wdata_oe_2x_r_8;
output 	wdp_wdata_oe_2x_r_9;
output 	wdp_wdata_oe_2x_r_10;
output 	wdp_wdata_oe_2x_r_11;
output 	wdp_wdata_oe_2x_r_12;
output 	wdp_wdata_oe_2x_r_13;
output 	wdp_wdata_oe_2x_r_14;
output 	wdp_wdata_oe_2x_r_15;
input 	control_wlat_r_0;
input 	control_doing_wr;
input 	Equal6;
input 	control_doing_wr1;
input 	control_doing_wr2;
output 	wd_lat_0;
output 	wd_lat_1;
output 	wd_lat_4;
output 	wd_lat_3;
output 	wd_lat_2;
input 	control_dqs_burst_0;
input 	dqs_burst_cas4;
input 	dqs_burst_cas3;
input 	GND_port;
input 	mem_clk_0;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altera_ddr_phy_alt_mem_phy altera_ddr_phy_alt_mem_phy_inst(
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.dm_ddio_dataout_0(dm_ddio_dataout_0),
	.dm_ddio_dataout_1(dm_ddio_dataout_1),
	.ddio_outa_0(ddio_outa_0),
	.ddio_outa_01(ddio_outa_01),
	.dq_ddio_dataout_0(dq_ddio_dataout_0),
	.dq_ddio_dataout_1(dq_ddio_dataout_1),
	.dq_ddio_dataout_2(dq_ddio_dataout_2),
	.dq_ddio_dataout_3(dq_ddio_dataout_3),
	.dq_ddio_dataout_4(dq_ddio_dataout_4),
	.dq_ddio_dataout_5(dq_ddio_dataout_5),
	.dq_ddio_dataout_6(dq_ddio_dataout_6),
	.dq_ddio_dataout_7(dq_ddio_dataout_7),
	.dq_ddio_dataout_8(dq_ddio_dataout_8),
	.dq_ddio_dataout_9(dq_ddio_dataout_9),
	.dq_ddio_dataout_10(dq_ddio_dataout_10),
	.dq_ddio_dataout_11(dq_ddio_dataout_11),
	.dq_ddio_dataout_12(dq_ddio_dataout_12),
	.dq_ddio_dataout_13(dq_ddio_dataout_13),
	.dq_ddio_dataout_14(dq_ddio_dataout_14),
	.dq_ddio_dataout_15(dq_ddio_dataout_15),
	.dqs_ddio_dataout_0(dqs_ddio_dataout_0),
	.wdp_wdqs_oe_2x_r_0(wdp_wdqs_oe_2x_r_0),
	.dqs_ddio_dataout_1(dqs_ddio_dataout_1),
	.wdp_wdqs_oe_2x_r_1(wdp_wdqs_oe_2x_r_1),
	.q_b_34(q_b_34),
	.q_b_32(q_b_32),
	.q_b_35(q_b_35),
	.q_b_33(q_b_33),
	.q_b_161(q_b_161),
	.q_b_01(q_b_01),
	.q_b_171(q_b_171),
	.q_b_110(q_b_110),
	.q_b_181(q_b_181),
	.q_b_210(q_b_210),
	.q_b_191(q_b_191),
	.q_b_36(q_b_36),
	.q_b_201(q_b_201),
	.q_b_41(q_b_41),
	.q_b_211(q_b_211),
	.q_b_51(q_b_51),
	.q_b_221(q_b_221),
	.q_b_61(q_b_61),
	.q_b_231(q_b_231),
	.q_b_71(q_b_71),
	.q_b_241(q_b_241),
	.q_b_81(q_b_81),
	.q_b_251(q_b_251),
	.q_b_91(q_b_91),
	.q_b_261(q_b_261),
	.q_b_101(q_b_101),
	.q_b_271(q_b_271),
	.q_b_111(q_b_111),
	.q_b_281(q_b_281),
	.q_b_121(q_b_121),
	.q_b_291(q_b_291),
	.q_b_131(q_b_131),
	.q_b_301(q_b_301),
	.q_b_141(q_b_141),
	.q_b_311(q_b_311),
	.q_b_151(q_b_151),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.reset_request_n(reset_request_n),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.control_doing_rd_0(control_doing_rd_0),
	.cs_n_0(cs_n_0),
	.a_0(a_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.ba_0(ba_0),
	.ba_1(ba_1),
	.ras_n(ras_n),
	.cas_n(cas_n),
	.we_n(we_n),
	.wdp_wdata_oe_2x_r_0(wdp_wdata_oe_2x_r_0),
	.wdp_wdata_oe_2x_r_1(wdp_wdata_oe_2x_r_1),
	.wdp_wdata_oe_2x_r_2(wdp_wdata_oe_2x_r_2),
	.wdp_wdata_oe_2x_r_3(wdp_wdata_oe_2x_r_3),
	.wdp_wdata_oe_2x_r_4(wdp_wdata_oe_2x_r_4),
	.wdp_wdata_oe_2x_r_5(wdp_wdata_oe_2x_r_5),
	.wdp_wdata_oe_2x_r_6(wdp_wdata_oe_2x_r_6),
	.wdp_wdata_oe_2x_r_7(wdp_wdata_oe_2x_r_7),
	.wdp_wdata_oe_2x_r_8(wdp_wdata_oe_2x_r_8),
	.wdp_wdata_oe_2x_r_9(wdp_wdata_oe_2x_r_9),
	.wdp_wdata_oe_2x_r_10(wdp_wdata_oe_2x_r_10),
	.wdp_wdata_oe_2x_r_11(wdp_wdata_oe_2x_r_11),
	.wdp_wdata_oe_2x_r_12(wdp_wdata_oe_2x_r_12),
	.wdp_wdata_oe_2x_r_13(wdp_wdata_oe_2x_r_13),
	.wdp_wdata_oe_2x_r_14(wdp_wdata_oe_2x_r_14),
	.wdp_wdata_oe_2x_r_15(wdp_wdata_oe_2x_r_15),
	.control_wlat_r_0(control_wlat_r_0),
	.control_doing_wr(control_doing_wr),
	.Equal6(Equal6),
	.control_doing_wr1(control_doing_wr1),
	.control_doing_wr2(control_doing_wr2),
	.wd_lat_0(wd_lat_0),
	.wd_lat_1(wd_lat_1),
	.wd_lat_4(wd_lat_4),
	.wd_lat_3(wd_lat_3),
	.wd_lat_2(wd_lat_2),
	.control_dqs_burst_0(control_dqs_burst_0),
	.dqs_burst_cas4(dqs_burst_cas4),
	.dqs_burst_cas3(dqs_burst_cas3),
	.GND_port(GND_port),
	.mem_clk_0(mem_clk_0),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy (
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dm_ddio_dataout_0,
	dm_ddio_dataout_1,
	ddio_outa_0,
	ddio_outa_01,
	dq_ddio_dataout_0,
	dq_ddio_dataout_1,
	dq_ddio_dataout_2,
	dq_ddio_dataout_3,
	dq_ddio_dataout_4,
	dq_ddio_dataout_5,
	dq_ddio_dataout_6,
	dq_ddio_dataout_7,
	dq_ddio_dataout_8,
	dq_ddio_dataout_9,
	dq_ddio_dataout_10,
	dq_ddio_dataout_11,
	dq_ddio_dataout_12,
	dq_ddio_dataout_13,
	dq_ddio_dataout_14,
	dq_ddio_dataout_15,
	dqs_ddio_dataout_0,
	wdp_wdqs_oe_2x_r_0,
	dqs_ddio_dataout_1,
	wdp_wdqs_oe_2x_r_1,
	q_b_34,
	q_b_32,
	q_b_35,
	q_b_33,
	q_b_161,
	q_b_01,
	q_b_171,
	q_b_110,
	q_b_181,
	q_b_210,
	q_b_191,
	q_b_36,
	q_b_201,
	q_b_41,
	q_b_211,
	q_b_51,
	q_b_221,
	q_b_61,
	q_b_231,
	q_b_71,
	q_b_241,
	q_b_81,
	q_b_251,
	q_b_91,
	q_b_261,
	q_b_101,
	q_b_271,
	q_b_111,
	q_b_281,
	q_b_121,
	q_b_291,
	q_b_131,
	q_b_301,
	q_b_141,
	q_b_311,
	q_b_151,
	seq_ac_add_1t_ac_lat_internal,
	ctl_rdata_valid_0,
	reset_request_n,
	ctl_init_success,
	reset_phy_clk_1x_n,
	control_doing_rd_0,
	cs_n_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	ba_0,
	ba_1,
	ras_n,
	cas_n,
	we_n,
	wdp_wdata_oe_2x_r_0,
	wdp_wdata_oe_2x_r_1,
	wdp_wdata_oe_2x_r_2,
	wdp_wdata_oe_2x_r_3,
	wdp_wdata_oe_2x_r_4,
	wdp_wdata_oe_2x_r_5,
	wdp_wdata_oe_2x_r_6,
	wdp_wdata_oe_2x_r_7,
	wdp_wdata_oe_2x_r_8,
	wdp_wdata_oe_2x_r_9,
	wdp_wdata_oe_2x_r_10,
	wdp_wdata_oe_2x_r_11,
	wdp_wdata_oe_2x_r_12,
	wdp_wdata_oe_2x_r_13,
	wdp_wdata_oe_2x_r_14,
	wdp_wdata_oe_2x_r_15,
	control_wlat_r_0,
	control_doing_wr,
	Equal6,
	control_doing_wr1,
	control_doing_wr2,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	control_dqs_burst_0,
	dqs_burst_cas4,
	dqs_burst_cas3,
	GND_port,
	mem_clk_0,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=1 */;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dm_ddio_dataout_0;
output 	dm_ddio_dataout_1;
output 	ddio_outa_0;
output 	ddio_outa_01;
output 	dq_ddio_dataout_0;
output 	dq_ddio_dataout_1;
output 	dq_ddio_dataout_2;
output 	dq_ddio_dataout_3;
output 	dq_ddio_dataout_4;
output 	dq_ddio_dataout_5;
output 	dq_ddio_dataout_6;
output 	dq_ddio_dataout_7;
output 	dq_ddio_dataout_8;
output 	dq_ddio_dataout_9;
output 	dq_ddio_dataout_10;
output 	dq_ddio_dataout_11;
output 	dq_ddio_dataout_12;
output 	dq_ddio_dataout_13;
output 	dq_ddio_dataout_14;
output 	dq_ddio_dataout_15;
output 	dqs_ddio_dataout_0;
output 	wdp_wdqs_oe_2x_r_0;
output 	dqs_ddio_dataout_1;
output 	wdp_wdqs_oe_2x_r_1;
input 	q_b_34;
input 	q_b_32;
input 	q_b_35;
input 	q_b_33;
input 	q_b_161;
input 	q_b_01;
input 	q_b_171;
input 	q_b_110;
input 	q_b_181;
input 	q_b_210;
input 	q_b_191;
input 	q_b_36;
input 	q_b_201;
input 	q_b_41;
input 	q_b_211;
input 	q_b_51;
input 	q_b_221;
input 	q_b_61;
input 	q_b_231;
input 	q_b_71;
input 	q_b_241;
input 	q_b_81;
input 	q_b_251;
input 	q_b_91;
input 	q_b_261;
input 	q_b_101;
input 	q_b_271;
input 	q_b_111;
input 	q_b_281;
input 	q_b_121;
input 	q_b_291;
input 	q_b_131;
input 	q_b_301;
input 	q_b_141;
input 	q_b_311;
input 	q_b_151;
output 	seq_ac_add_1t_ac_lat_internal;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	ctl_init_success;
output 	reset_phy_clk_1x_n;
input 	control_doing_rd_0;
input 	cs_n_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	ba_0;
input 	ba_1;
input 	ras_n;
input 	cas_n;
input 	we_n;
output 	wdp_wdata_oe_2x_r_0;
output 	wdp_wdata_oe_2x_r_1;
output 	wdp_wdata_oe_2x_r_2;
output 	wdp_wdata_oe_2x_r_3;
output 	wdp_wdata_oe_2x_r_4;
output 	wdp_wdata_oe_2x_r_5;
output 	wdp_wdata_oe_2x_r_6;
output 	wdp_wdata_oe_2x_r_7;
output 	wdp_wdata_oe_2x_r_8;
output 	wdp_wdata_oe_2x_r_9;
output 	wdp_wdata_oe_2x_r_10;
output 	wdp_wdata_oe_2x_r_11;
output 	wdp_wdata_oe_2x_r_12;
output 	wdp_wdata_oe_2x_r_13;
output 	wdp_wdata_oe_2x_r_14;
output 	wdp_wdata_oe_2x_r_15;
input 	control_wlat_r_0;
input 	control_doing_wr;
input 	Equal6;
input 	control_doing_wr1;
input 	control_doing_wr2;
output 	wd_lat_0;
output 	wd_lat_1;
output 	wd_lat_4;
output 	wd_lat_3;
output 	wd_lat_2;
input 	control_dqs_burst_0;
input 	dqs_burst_cas4;
input 	dqs_burst_cas3;
input 	GND_port;
input 	mem_clk_0;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \clk|pll|altpll_component|auto_generated|clk[2] ;
wire \clk|pll|altpll_component|auto_generated|clk[3] ;
wire \clk|pll|altpll_component|auto_generated|clk[4] ;
wire \seq_wrapper|seq_inst|seq_ac_addr[2]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[3]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[4]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[5]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[8]~q ;
wire \rdv_pipe|rd_addr[0]~q ;
wire \rdp|rd_ram_rd_addr[1]~q ;
wire \rdp|rd_ram_rd_addr[2]~q ;
wire \rdp|rd_ram_rd_addr[3]~q ;
wire \clk|ac_clk_pipe_2x|ams_pipe[1]~q ;
wire \seq_wrapper|seq_inst|ctrl|ctl_init_success~q ;
wire \full_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q ;
wire \full_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q ;
wire \full_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ;
wire \full_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ;
wire \clk|resync_clk_pipe|ams_pipe[1]~q ;
wire \seq_wrapper|seq_inst|seq_rdv_doing_rd[0]~q ;
wire \seq_wrapper|seq_inst|seq_rdv_doing_rd[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_cke[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[8]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[10]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ras_n[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_cas_n[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_we_n[0]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ;
wire \seq_wrapper|seq_inst|seq_wdp_ovride~2_combout ;
wire \dpio|dio_rdata_h_2x[0]~q ;
wire \dpio|dio_rdata_h_2x[1]~q ;
wire \dpio|dio_rdata_h_2x[2]~q ;
wire \dpio|dio_rdata_h_2x[3]~q ;
wire \dpio|dio_rdata_h_2x[4]~q ;
wire \dpio|dio_rdata_h_2x[5]~q ;
wire \dpio|dio_rdata_h_2x[6]~q ;
wire \dpio|dio_rdata_h_2x[7]~q ;
wire \dpio|dio_rdata_h_2x[8]~q ;
wire \dpio|dio_rdata_h_2x[9]~q ;
wire \dpio|dio_rdata_h_2x[10]~q ;
wire \dpio|dio_rdata_h_2x[11]~q ;
wire \dpio|dio_rdata_h_2x[12]~q ;
wire \dpio|dio_rdata_h_2x[13]~q ;
wire \dpio|dio_rdata_h_2x[14]~q ;
wire \dpio|dio_rdata_h_2x[15]~q ;
wire \dpio|dio_rdata_l_2x[0]~q ;
wire \dpio|dio_rdata_l_2x[1]~q ;
wire \dpio|dio_rdata_l_2x[2]~q ;
wire \dpio|dio_rdata_l_2x[3]~q ;
wire \dpio|dio_rdata_l_2x[4]~q ;
wire \dpio|dio_rdata_l_2x[5]~q ;
wire \dpio|dio_rdata_l_2x[6]~q ;
wire \dpio|dio_rdata_l_2x[7]~q ;
wire \dpio|dio_rdata_l_2x[8]~q ;
wire \dpio|dio_rdata_l_2x[9]~q ;
wire \dpio|dio_rdata_l_2x[10]~q ;
wire \dpio|dio_rdata_l_2x[11]~q ;
wire \dpio|dio_rdata_l_2x[12]~q ;
wire \dpio|dio_rdata_l_2x[13]~q ;
wire \dpio|dio_rdata_l_2x[14]~q ;
wire \dpio|dio_rdata_l_2x[15]~q ;
wire \seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ;
wire \rdp|Add2~0_combout ;
wire \seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ;
wire \seq_wrapper|seq_inst|seq_pll_start_reconfig~q ;
wire \seq_wrapper|seq_inst|seq_mem_clk_disable~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q ;
wire \full_rate_wdp_gen.wdp|dq_oe_2x[0]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ;
wire \full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ;
wire \full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ;
wire \full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdqs_2x[1]~q ;
wire \full_rate_wdp_gen.wdp|wdp_wdqs_oe_2x[0]~q ;
wire \seq_wrapper|seq_inst|seq_pll_select[2]~q ;
wire \seq_wrapper|seq_inst|seq_pll_select[0]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[9]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[10]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[11]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[12]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[13]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[14]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[15]~q ;
wire \rdv_pipe|seq_rdata_valid[0]~q ;
wire \clk|phs_shft_busy~q ;
wire \mmc|mimic_done_out~q ;
wire \clk|measure_clk_pipe|ams_pipe[1]~q ;
wire \seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ;
wire \mmc|mimic_value_captured~q ;
wire \clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|input_cell_h[0]~q ;


altera_ddr_altera_ddr_phy_alt_mem_phy_rdata_valid rdv_pipe(
	.clk_1(clk_1),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rd_addr_0(\rdv_pipe|rd_addr[0]~q ),
	.rd_ram_rd_addr_1(\rdp|rd_ram_rd_addr[1]~q ),
	.rd_ram_rd_addr_2(\rdp|rd_ram_rd_addr[2]~q ),
	.rd_ram_rd_addr_3(\rdp|rd_ram_rd_addr[3]~q ),
	.seq_rdv_doing_rd_0(\seq_wrapper|seq_inst|seq_rdv_doing_rd[0]~q ),
	.seq_rdv_doing_rd_1(\seq_wrapper|seq_inst|seq_rdv_doing_rd[1]~q ),
	.control_doing_rd_0(control_doing_rd_0),
	.seq_rdata_valid_lat_dec(\seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ),
	.Add2(\rdp|Add2~0_combout ),
	.seq_rdata_valid_0(\rdv_pipe|seq_rdata_valid[0]~q ));

altera_ddr_altera_ddr_phy_alt_mem_phy_clk_reset clk(
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_2(\clk|pll|altpll_component|auto_generated|clk[2] ),
	.clk_3(\clk|pll|altpll_component|auto_generated|clk[3] ),
	.clk_4(\clk|pll|altpll_component|auto_generated|clk[4] ),
	.ddio_outa_0(ddio_outa_0),
	.ddio_outa_01(ddio_outa_01),
	.reset_request_n(reset_request_n),
	.reset_phy_clk_1x_n1(reset_phy_clk_1x_n),
	.ams_pipe_1(\clk|ac_clk_pipe_2x|ams_pipe[1]~q ),
	.ams_pipe_11(\clk|resync_clk_pipe|ams_pipe[1]~q ),
	.seq_pll_inc_dec_n(\seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig(\seq_wrapper|seq_inst|seq_pll_start_reconfig~q ),
	.seq_mem_clk_disable(\seq_wrapper|seq_inst|seq_mem_clk_disable~q ),
	.seq_pll_select({\seq_wrapper|seq_inst|seq_pll_select[2]~q ,gnd,\seq_wrapper|seq_inst|seq_pll_select[0]~q }),
	.phs_shft_busy1(\clk|phs_shft_busy~q ),
	.ams_pipe_12(\clk|measure_clk_pipe|ams_pipe[1]~q ),
	.input_cell_h_0(\clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|input_cell_h[0]~q ),
	.mem_clk_0(mem_clk_0),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

altera_ddr_altera_ddr_phy_alt_mem_phy_mimic mmc(
	.measure_clk(\clk|pll|altpll_component|auto_generated|clk[4] ),
	.mimic_done_out1(\mmc|mimic_done_out~q ),
	.reset_measure_clk_n(\clk|measure_clk_pipe|ams_pipe[1]~q ),
	.seq_mmc_start(\seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ),
	.mimic_value_captured1(\mmc|mimic_value_captured~q ),
	.mimic_data_in(\clk|DDR_CLK_OUT[0].ddr_clk_out_p|auto_generated|input_cell_h[0]~q ));

altera_ddr_altera_ddr_phy_alt_mem_phy_seq_wrapper seq_wrapper(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk_1(clk_1),
	.seq_ac_addr_2(\seq_wrapper|seq_inst|seq_ac_addr[2]~q ),
	.seq_ac_addr_3(\seq_wrapper|seq_inst|seq_ac_addr[3]~q ),
	.seq_ac_addr_4(\seq_wrapper|seq_inst|seq_ac_addr[4]~q ),
	.seq_ac_addr_5(\seq_wrapper|seq_inst|seq_ac_addr[5]~q ),
	.dgwb_wdata_24(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ),
	.dgwb_wdata_8(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[8]~q ),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.ctl_init_success1(\seq_wrapper|seq_inst|ctrl|ctl_init_success~q ),
	.seq_rdv_doing_rd_0(\seq_wrapper|seq_inst|seq_rdv_doing_rd[0]~q ),
	.seq_rdv_doing_rd_1(\seq_wrapper|seq_inst|seq_rdv_doing_rd[1]~q ),
	.seq_ac_cs_n_0(\seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ),
	.seq_ac_cke_0(\seq_wrapper|seq_inst|seq_ac_cke[0]~q ),
	.seq_ac_addr_0(\seq_wrapper|seq_inst|seq_ac_addr[0]~q ),
	.seq_ac_addr_1(\seq_wrapper|seq_inst|seq_ac_addr[1]~q ),
	.seq_ac_addr_8(\seq_wrapper|seq_inst|seq_ac_addr[8]~q ),
	.seq_ac_addr_10(\seq_wrapper|seq_inst|seq_ac_addr[10]~q ),
	.seq_ac_ba_0(\seq_wrapper|seq_inst|seq_ac_ba[0]~q ),
	.seq_ac_ba_1(\seq_wrapper|seq_inst|seq_ac_ba[1]~q ),
	.seq_ac_ras_n_0(\seq_wrapper|seq_inst|seq_ac_ras_n[0]~q ),
	.seq_ac_cas_n_0(\seq_wrapper|seq_inst|seq_ac_cas_n[0]~q ),
	.seq_ac_we_n_0(\seq_wrapper|seq_inst|seq_ac_we_n[0]~q ),
	.dgwb_wdp_ovride(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ),
	.seq_wdp_ovride(\seq_wrapper|seq_inst|seq_wdp_ovride~2_combout ),
	.seq_rdata_valid_lat_dec(\seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ),
	.seq_pll_inc_dec_n(\seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig(\seq_wrapper|seq_inst|seq_pll_start_reconfig~q ),
	.seq_mem_clk_disable(\seq_wrapper|seq_inst|seq_mem_clk_disable~q ),
	.wd_lat_0(wd_lat_0),
	.wd_lat_1(wd_lat_1),
	.wd_lat_4(wd_lat_4),
	.wd_lat_3(wd_lat_3),
	.wd_lat_2(wd_lat_2),
	.seq_pll_select_2(\seq_wrapper|seq_inst|seq_pll_select[2]~q ),
	.seq_pll_select_0(\seq_wrapper|seq_inst|seq_pll_select[0]~q ),
	.dgwb_wdata_25(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ),
	.dgwb_wdata_9(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[9]~q ),
	.dgwb_wdata_26(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ),
	.dgwb_wdata_10(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[10]~q ),
	.dgwb_wdata_27(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ),
	.dgwb_wdata_11(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[11]~q ),
	.dgwb_wdata_28(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ),
	.dgwb_wdata_12(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[12]~q ),
	.dgwb_wdata_29(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ),
	.dgwb_wdata_13(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[13]~q ),
	.dgwb_wdata_30(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ),
	.dgwb_wdata_14(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[14]~q ),
	.dgwb_wdata_31(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ),
	.dgwb_wdata_15(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[15]~q ),
	.seq_rdata_valid_0(\rdv_pipe|seq_rdata_valid[0]~q ),
	.phs_shft_busy(\clk|phs_shft_busy~q ),
	.mimic_done_out(\mmc|mimic_done_out~q ),
	.seq_mmc_start(\seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ),
	.mimic_value_captured(\mmc|mimic_value_captured~q ),
	.GND_port(GND_port));

altera_ddr_altera_ddr_phy_alt_mem_phy_read_dp rdp(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk_1(clk_1),
	.clk_3(\clk|pll|altpll_component|auto_generated|clk[3] ),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rd_addr_0(\rdv_pipe|rd_addr[0]~q ),
	.rd_ram_rd_addr_1(\rdp|rd_ram_rd_addr[1]~q ),
	.rd_ram_rd_addr_2(\rdp|rd_ram_rd_addr[2]~q ),
	.rd_ram_rd_addr_3(\rdp|rd_ram_rd_addr[3]~q ),
	.reset_resync_clk_2x_n(\clk|resync_clk_pipe|ams_pipe[1]~q ),
	.dio_rdata_h_2x({\dpio|dio_rdata_h_2x[15]~q ,\dpio|dio_rdata_h_2x[14]~q ,\dpio|dio_rdata_h_2x[13]~q ,\dpio|dio_rdata_h_2x[12]~q ,\dpio|dio_rdata_h_2x[11]~q ,\dpio|dio_rdata_h_2x[10]~q ,\dpio|dio_rdata_h_2x[9]~q ,\dpio|dio_rdata_h_2x[8]~q ,\dpio|dio_rdata_h_2x[7]~q ,
\dpio|dio_rdata_h_2x[6]~q ,\dpio|dio_rdata_h_2x[5]~q ,\dpio|dio_rdata_h_2x[4]~q ,\dpio|dio_rdata_h_2x[3]~q ,\dpio|dio_rdata_h_2x[2]~q ,\dpio|dio_rdata_h_2x[1]~q ,\dpio|dio_rdata_h_2x[0]~q }),
	.dio_rdata_l_2x({\dpio|dio_rdata_l_2x[15]~q ,\dpio|dio_rdata_l_2x[14]~q ,\dpio|dio_rdata_l_2x[13]~q ,\dpio|dio_rdata_l_2x[12]~q ,\dpio|dio_rdata_l_2x[11]~q ,\dpio|dio_rdata_l_2x[10]~q ,\dpio|dio_rdata_l_2x[9]~q ,\dpio|dio_rdata_l_2x[8]~q ,\dpio|dio_rdata_l_2x[7]~q ,
\dpio|dio_rdata_l_2x[6]~q ,\dpio|dio_rdata_l_2x[5]~q ,\dpio|dio_rdata_l_2x[4]~q ,\dpio|dio_rdata_l_2x[3]~q ,\dpio|dio_rdata_l_2x[2]~q ,\dpio|dio_rdata_l_2x[1]~q ,\dpio|dio_rdata_l_2x[0]~q }),
	.Add2(\rdp|Add2~0_combout ));

altera_ddr_altera_ddr_phy_alt_mem_phy_write_dp_fr \full_rate_wdp_gen.wdp (
	.phy_clk_1x(clk_1),
	.q_b_34(q_b_34),
	.q_b_32(q_b_32),
	.q_b_35(q_b_35),
	.q_b_33(q_b_33),
	.q_b_16(q_b_161),
	.dgwb_wdata_24(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ),
	.q_b_0(q_b_01),
	.dgwb_wdata_8(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[8]~q ),
	.q_b_17(q_b_171),
	.q_b_1(q_b_110),
	.q_b_18(q_b_181),
	.q_b_2(q_b_210),
	.q_b_19(q_b_191),
	.q_b_3(q_b_36),
	.q_b_20(q_b_201),
	.q_b_4(q_b_41),
	.q_b_21(q_b_211),
	.q_b_5(q_b_51),
	.q_b_22(q_b_221),
	.q_b_6(q_b_61),
	.q_b_23(q_b_231),
	.q_b_7(q_b_71),
	.q_b_24(q_b_241),
	.q_b_8(q_b_81),
	.q_b_25(q_b_251),
	.q_b_9(q_b_91),
	.q_b_26(q_b_261),
	.q_b_10(q_b_101),
	.q_b_27(q_b_271),
	.q_b_11(q_b_111),
	.q_b_28(q_b_281),
	.q_b_12(q_b_121),
	.q_b_29(q_b_291),
	.q_b_13(q_b_131),
	.q_b_30(q_b_301),
	.q_b_14(q_b_141),
	.q_b_31(q_b_311),
	.q_b_15(q_b_151),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.ctl_init_success(\seq_wrapper|seq_inst|ctrl|ctl_init_success~q ),
	.wdp_dm_l_2x_0(\full_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q ),
	.wdp_dm_h_2x_0(\full_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q ),
	.wdp_dm_l_2x_1(\full_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ),
	.wdp_dm_h_2x_1(\full_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ),
	.control_wlat_r_0(control_wlat_r_0),
	.control_doing_wr(control_doing_wr),
	.Equal6(Equal6),
	.control_doing_wr1(control_doing_wr1),
	.control_doing_wr2(control_doing_wr2),
	.dgwb_wdp_ovride(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ),
	.seq_wdp_ovride(\seq_wrapper|seq_inst|seq_wdp_ovride~2_combout ),
	.wdp_wdata_l_2x_0(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q ),
	.wdp_wdata_h_2x_0(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q ),
	.dq_oe_2x_0(\full_rate_wdp_gen.wdp|dq_oe_2x[0]~q ),
	.wdp_wdata_l_2x_1(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ),
	.wdp_wdata_h_2x_1(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ),
	.wdp_wdata_l_2x_2(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ),
	.wdp_wdata_h_2x_2(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ),
	.wdp_wdata_l_2x_3(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ),
	.wdp_wdata_h_2x_3(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ),
	.wdp_wdata_l_2x_4(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ),
	.wdp_wdata_h_2x_4(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ),
	.dq_oe_2x_1(\full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ),
	.wdp_wdata_l_2x_5(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ),
	.wdp_wdata_h_2x_5(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ),
	.wdp_wdata_l_2x_6(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ),
	.wdp_wdata_h_2x_6(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ),
	.wdp_wdata_l_2x_7(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ),
	.wdp_wdata_h_2x_7(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ),
	.wdp_wdata_l_2x_8(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ),
	.wdp_wdata_h_2x_8(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ),
	.dq_oe_2x_2(\full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ),
	.wdp_wdata_l_2x_9(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ),
	.wdp_wdata_h_2x_9(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ),
	.wdp_wdata_l_2x_10(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ),
	.wdp_wdata_h_2x_10(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ),
	.wdp_wdata_l_2x_11(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ),
	.wdp_wdata_h_2x_11(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ),
	.wdp_wdata_l_2x_12(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ),
	.wdp_wdata_h_2x_12(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ),
	.dq_oe_2x_3(\full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ),
	.wdp_wdata_l_2x_13(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ),
	.wdp_wdata_h_2x_13(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ),
	.wdp_wdata_l_2x_14(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ),
	.wdp_wdata_h_2x_14(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ),
	.wdp_wdata_l_2x_15(\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ),
	.wdp_wdata_h_2x_15(\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ),
	.wdp_wdqs_2x_1(\full_rate_wdp_gen.wdp|wdp_wdqs_2x[1]~q ),
	.wdp_wdqs_oe_2x_0(\full_rate_wdp_gen.wdp|wdp_wdqs_oe_2x[0]~q ),
	.dgwb_wdata_25(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ),
	.dgwb_wdata_9(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[9]~q ),
	.dgwb_wdata_26(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ),
	.dgwb_wdata_10(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[10]~q ),
	.dgwb_wdata_27(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ),
	.dgwb_wdata_11(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[11]~q ),
	.dgwb_wdata_28(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ),
	.dgwb_wdata_12(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[12]~q ),
	.dgwb_wdata_29(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ),
	.dgwb_wdata_13(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[13]~q ),
	.dgwb_wdata_30(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ),
	.dgwb_wdata_14(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[14]~q ),
	.dgwb_wdata_31(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ),
	.dgwb_wdata_15(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[15]~q ),
	.control_dqs_burst_0(control_dqs_burst_0),
	.dqs_burst_cas4(dqs_burst_cas4),
	.dqs_burst_cas3(dqs_burst_cas3));

altera_ddr_altera_ddr_phy_alt_mem_phy_addr_cmd \full_rate_adc_gen.adc (
	.clk_1(clk_1),
	.clk_2(\clk|pll|altpll_component|auto_generated|clk[2] ),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.seq_ac_addr_2(\seq_wrapper|seq_inst|seq_ac_addr[2]~q ),
	.seq_ac_addr_3(\seq_wrapper|seq_inst|seq_ac_addr[3]~q ),
	.seq_ac_addr_4(\seq_wrapper|seq_inst|seq_ac_addr[4]~q ),
	.seq_ac_addr_5(\seq_wrapper|seq_inst|seq_ac_addr[5]~q ),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.ams_pipe_1(\clk|ac_clk_pipe_2x|ams_pipe[1]~q ),
	.seq_ac_cs_n_0(\seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ),
	.cs_n_0(cs_n_0),
	.seq_ac_cke_0(\seq_wrapper|seq_inst|seq_ac_cke[0]~q ),
	.a_0(a_0),
	.seq_ac_addr_0(\seq_wrapper|seq_inst|seq_ac_addr[0]~q ),
	.a_1(a_1),
	.seq_ac_addr_1(\seq_wrapper|seq_inst|seq_ac_addr[1]~q ),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.seq_ac_addr_8(\seq_wrapper|seq_inst|seq_ac_addr[8]~q ),
	.a_9(a_9),
	.a_10(a_10),
	.seq_ac_addr_10(\seq_wrapper|seq_inst|seq_ac_addr[10]~q ),
	.a_11(a_11),
	.a_12(a_12),
	.seq_ac_ba_0(\seq_wrapper|seq_inst|seq_ac_ba[0]~q ),
	.ba_0(ba_0),
	.seq_ac_ba_1(\seq_wrapper|seq_inst|seq_ac_ba[1]~q ),
	.ba_1(ba_1),
	.seq_ac_ras_n_0(\seq_wrapper|seq_inst|seq_ac_ras_n[0]~q ),
	.ras_n(ras_n),
	.seq_ac_cas_n_0(\seq_wrapper|seq_inst|seq_ac_cas_n[0]~q ),
	.cas_n(cas_n),
	.seq_ac_we_n_0(\seq_wrapper|seq_inst|seq_ac_we_n[0]~q ),
	.we_n(we_n));

altera_ddr_altera_ddr_phy_alt_mem_phy_dp_io dpio(
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.mem_clk_2x(clk_1),
	.write_clk_2x(\clk|pll|altpll_component|auto_generated|clk[2] ),
	.clk_3(\clk|pll|altpll_component|auto_generated|clk[3] ),
	.dm_ddio_dataout_0(dm_ddio_dataout_0),
	.dm_ddio_dataout_1(dm_ddio_dataout_1),
	.dq_ddio_dataout_0(dq_ddio_dataout_0),
	.dq_ddio_dataout_1(dq_ddio_dataout_1),
	.dq_ddio_dataout_2(dq_ddio_dataout_2),
	.dq_ddio_dataout_3(dq_ddio_dataout_3),
	.dq_ddio_dataout_4(dq_ddio_dataout_4),
	.dq_ddio_dataout_5(dq_ddio_dataout_5),
	.dq_ddio_dataout_6(dq_ddio_dataout_6),
	.dq_ddio_dataout_7(dq_ddio_dataout_7),
	.dq_ddio_dataout_8(dq_ddio_dataout_8),
	.dq_ddio_dataout_9(dq_ddio_dataout_9),
	.dq_ddio_dataout_10(dq_ddio_dataout_10),
	.dq_ddio_dataout_11(dq_ddio_dataout_11),
	.dq_ddio_dataout_12(dq_ddio_dataout_12),
	.dq_ddio_dataout_13(dq_ddio_dataout_13),
	.dq_ddio_dataout_14(dq_ddio_dataout_14),
	.dq_ddio_dataout_15(dq_ddio_dataout_15),
	.dqs_ddio_dataout_0(dqs_ddio_dataout_0),
	.wdp_wdqs_oe_2x_r_0(wdp_wdqs_oe_2x_r_0),
	.dqs_ddio_dataout_1(dqs_ddio_dataout_1),
	.wdp_wdqs_oe_2x_r_1(wdp_wdqs_oe_2x_r_1),
	.wdp_dm_l_2x({\full_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ,\full_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q }),
	.wdp_dm_h_2x({\full_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ,\full_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q }),
	.ams_pipe_1(\clk|resync_clk_pipe|ams_pipe[1]~q ),
	.wdp_wdata_oe_2x_r_0(wdp_wdata_oe_2x_r_0),
	.wdp_wdata_oe_2x_r_1(wdp_wdata_oe_2x_r_1),
	.wdp_wdata_oe_2x_r_2(wdp_wdata_oe_2x_r_2),
	.wdp_wdata_oe_2x_r_3(wdp_wdata_oe_2x_r_3),
	.wdp_wdata_oe_2x_r_4(wdp_wdata_oe_2x_r_4),
	.wdp_wdata_oe_2x_r_5(wdp_wdata_oe_2x_r_5),
	.wdp_wdata_oe_2x_r_6(wdp_wdata_oe_2x_r_6),
	.wdp_wdata_oe_2x_r_7(wdp_wdata_oe_2x_r_7),
	.wdp_wdata_oe_2x_r_8(wdp_wdata_oe_2x_r_8),
	.wdp_wdata_oe_2x_r_9(wdp_wdata_oe_2x_r_9),
	.wdp_wdata_oe_2x_r_10(wdp_wdata_oe_2x_r_10),
	.wdp_wdata_oe_2x_r_11(wdp_wdata_oe_2x_r_11),
	.wdp_wdata_oe_2x_r_12(wdp_wdata_oe_2x_r_12),
	.wdp_wdata_oe_2x_r_13(wdp_wdata_oe_2x_r_13),
	.wdp_wdata_oe_2x_r_14(wdp_wdata_oe_2x_r_14),
	.wdp_wdata_oe_2x_r_15(wdp_wdata_oe_2x_r_15),
	.dio_rdata_h_2x_0(\dpio|dio_rdata_h_2x[0]~q ),
	.dio_rdata_h_2x_1(\dpio|dio_rdata_h_2x[1]~q ),
	.dio_rdata_h_2x_2(\dpio|dio_rdata_h_2x[2]~q ),
	.dio_rdata_h_2x_3(\dpio|dio_rdata_h_2x[3]~q ),
	.dio_rdata_h_2x_4(\dpio|dio_rdata_h_2x[4]~q ),
	.dio_rdata_h_2x_5(\dpio|dio_rdata_h_2x[5]~q ),
	.dio_rdata_h_2x_6(\dpio|dio_rdata_h_2x[6]~q ),
	.dio_rdata_h_2x_7(\dpio|dio_rdata_h_2x[7]~q ),
	.dio_rdata_h_2x_8(\dpio|dio_rdata_h_2x[8]~q ),
	.dio_rdata_h_2x_9(\dpio|dio_rdata_h_2x[9]~q ),
	.dio_rdata_h_2x_10(\dpio|dio_rdata_h_2x[10]~q ),
	.dio_rdata_h_2x_11(\dpio|dio_rdata_h_2x[11]~q ),
	.dio_rdata_h_2x_12(\dpio|dio_rdata_h_2x[12]~q ),
	.dio_rdata_h_2x_13(\dpio|dio_rdata_h_2x[13]~q ),
	.dio_rdata_h_2x_14(\dpio|dio_rdata_h_2x[14]~q ),
	.dio_rdata_h_2x_15(\dpio|dio_rdata_h_2x[15]~q ),
	.dio_rdata_l_2x_0(\dpio|dio_rdata_l_2x[0]~q ),
	.dio_rdata_l_2x_1(\dpio|dio_rdata_l_2x[1]~q ),
	.dio_rdata_l_2x_2(\dpio|dio_rdata_l_2x[2]~q ),
	.dio_rdata_l_2x_3(\dpio|dio_rdata_l_2x[3]~q ),
	.dio_rdata_l_2x_4(\dpio|dio_rdata_l_2x[4]~q ),
	.dio_rdata_l_2x_5(\dpio|dio_rdata_l_2x[5]~q ),
	.dio_rdata_l_2x_6(\dpio|dio_rdata_l_2x[6]~q ),
	.dio_rdata_l_2x_7(\dpio|dio_rdata_l_2x[7]~q ),
	.dio_rdata_l_2x_8(\dpio|dio_rdata_l_2x[8]~q ),
	.dio_rdata_l_2x_9(\dpio|dio_rdata_l_2x[9]~q ),
	.dio_rdata_l_2x_10(\dpio|dio_rdata_l_2x[10]~q ),
	.dio_rdata_l_2x_11(\dpio|dio_rdata_l_2x[11]~q ),
	.dio_rdata_l_2x_12(\dpio|dio_rdata_l_2x[12]~q ),
	.dio_rdata_l_2x_13(\dpio|dio_rdata_l_2x[13]~q ),
	.dio_rdata_l_2x_14(\dpio|dio_rdata_l_2x[14]~q ),
	.dio_rdata_l_2x_15(\dpio|dio_rdata_l_2x[15]~q ),
	.wdp_wdata_l_2x({\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q }),
	.wdp_wdata_h_2x({\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ,\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ,
\full_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q }),
	.wdp_wdata_oe_2x({\full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[3]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ,
\full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[2]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[1]~q ,
\full_rate_wdp_gen.wdp|dq_oe_2x[0]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[0]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[0]~q ,\full_rate_wdp_gen.wdp|dq_oe_2x[0]~q }),
	.wdp_wdqs_2x({\full_rate_wdp_gen.wdp|wdp_wdqs_2x[1]~q ,\full_rate_wdp_gen.wdp|wdp_wdqs_2x[1]~q }),
	.wdp_wdqs_oe_2x({\full_rate_wdp_gen.wdp|wdp_wdqs_oe_2x[0]~q ,\full_rate_wdp_gen.wdp|wdp_wdqs_oe_2x[0]~q }));

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_addr_cmd (
	clk_1,
	clk_2,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	seq_ac_addr_2,
	seq_ac_addr_3,
	seq_ac_addr_4,
	seq_ac_addr_5,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	ams_pipe_1,
	seq_ac_cs_n_0,
	cs_n_0,
	seq_ac_cke_0,
	a_0,
	seq_ac_addr_0,
	a_1,
	seq_ac_addr_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	seq_ac_addr_8,
	a_9,
	a_10,
	seq_ac_addr_10,
	a_11,
	a_12,
	seq_ac_ba_0,
	ba_0,
	seq_ac_ba_1,
	ba_1,
	seq_ac_ras_n_0,
	ras_n,
	seq_ac_cas_n_0,
	cas_n,
	seq_ac_we_n_0,
	we_n)/* synthesis synthesis_greybox=1 */;
input 	clk_1;
input 	clk_2;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
input 	seq_ac_addr_2;
input 	seq_ac_addr_3;
input 	seq_ac_addr_4;
input 	seq_ac_addr_5;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	ams_pipe_1;
input 	seq_ac_cs_n_0;
input 	cs_n_0;
input 	seq_ac_cke_0;
input 	a_0;
input 	seq_ac_addr_0;
input 	a_1;
input 	seq_ac_addr_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	seq_ac_addr_8;
input 	a_9;
input 	a_10;
input 	seq_ac_addr_10;
input 	a_11;
input 	a_12;
input 	seq_ac_ba_0;
input 	ba_0;
input 	seq_ac_ba_1;
input 	ba_1;
input 	seq_ac_ras_n_0;
input 	ras_n;
input 	seq_ac_cas_n_0;
input 	cas_n;
input 	seq_ac_we_n_0;
input 	we_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altera_ddr_phy_alt_mem_phy_ac_17 \cs_n[0].cs_n_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_0),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.ams_pipe_1(ams_pipe_1),
	.seq_ac_cs_n_0(seq_ac_cs_n_0),
	.cs_n_0(cs_n_0));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_18 ras_n_struct(
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_017),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_ras_n_0(seq_ac_ras_n_0),
	.ras_n(ras_n));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_19 we_n_struct(
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_019),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_we_n_0(seq_ac_we_n_0),
	.we_n(we_n));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac \addr[0].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_02),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_0(a_0),
	.seq_ac_addr_0(seq_ac_addr_0));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_4 \addr[1].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_03),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_1(a_1),
	.seq_ac_addr_1(seq_ac_addr_1));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_5 \addr[2].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_04),
	.seq_ac_addr_2(seq_ac_addr_2),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_2(a_2));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_6 \addr[3].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_05),
	.seq_ac_addr_3(seq_ac_addr_3),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_3(a_3));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_7 \addr[4].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_06),
	.seq_ac_addr_4(seq_ac_addr_4),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_4(a_4));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_8 \addr[5].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_07),
	.seq_ac_addr_5(seq_ac_addr_5),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_5(a_5));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_9 \addr[6].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_08),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_addr_0(seq_ac_addr_0),
	.a_6(a_6));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_10 \addr[7].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_09),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_addr_0(seq_ac_addr_0),
	.a_7(a_7));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_11 \addr[8].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_010),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_8(a_8),
	.seq_ac_addr_8(seq_ac_addr_8));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_12 \addr[9].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_011),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_addr_0(seq_ac_addr_0),
	.a_9(a_9));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_1 \addr[10].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_012),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.a_10(a_10),
	.seq_ac_addr_10(seq_ac_addr_10));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_2 \addr[11].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_013),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_addr_0(seq_ac_addr_0),
	.a_11(a_11));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_3 \addr[12].addr_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_014),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_addr_0(seq_ac_addr_0),
	.a_12(a_12));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_13 \ba[0].ba_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_015),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_ba_0(seq_ac_ba_0),
	.ba_0(ba_0));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_14 \ba[1].ba_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_016),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_ba_1(seq_ac_ba_1),
	.ba_1(ba_1));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_15 cas_n_struct(
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_018),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.seq_ac_cas_n_0(seq_ac_cas_n_0),
	.cas_n(cas_n));

altera_ddr_altera_ddr_phy_alt_mem_phy_ac_16 \cke[0].cke_struct (
	.phy_clk_1x(clk_1),
	.clk_2(clk_2),
	.dataout_0(dataout_01),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success(ctl_init_success),
	.ams_pipe_1(ams_pipe_1),
	.seq_ac_cke_0(seq_ac_cke_0));

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_0,
	seq_ac_addr_0)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_0;
input 	seq_ac_addr_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_1 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_0),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_1 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_10,
	seq_ac_addr_10)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_10;
input 	seq_ac_addr_10;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_2 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_10),
	.datab(seq_ac_addr_10),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_2 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_1 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_2 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_addr_0,
	a_11)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_addr_0;
input 	a_11;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_3 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_11),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_3 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_2 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_2 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_3 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_addr_0,
	a_12)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_addr_0;
input 	a_12;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_4 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_12),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_4 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_3 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_3 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_4 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_1,
	seq_ac_addr_1)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_1;
input 	seq_ac_addr_1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_5 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_1),
	.datab(seq_ac_addr_1),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_5 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_4 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_4 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_5 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_addr_2,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_2)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_addr_2;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_2;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_6 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_2),
	.datab(seq_ac_addr_2),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_6 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_5 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_5 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_6 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_addr_3,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_3)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_addr_3;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_3;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_7 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_3),
	.datab(seq_ac_addr_3),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_7 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_6 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_6 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_7 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_addr_4,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_4)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_addr_4;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_4;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_8 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_4),
	.datab(seq_ac_addr_4),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_8 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_7 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_7 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_8 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_addr_5,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_5)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_addr_5;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_5;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_9 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_5),
	.datab(seq_ac_addr_5),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_9 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_8 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_8 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_9 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_addr_0,
	a_6)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_addr_0;
input 	a_6;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_10 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_6),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_10 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_9 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_9 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_10 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_addr_0,
	a_7)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_addr_0;
input 	a_7;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_11 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_7),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_11 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_10 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_10 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_11 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	a_8,
	seq_ac_addr_8)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	a_8;
input 	seq_ac_addr_8;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_12 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_8),
	.datab(seq_ac_addr_8),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_12 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_11 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_11 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_12 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_addr_0,
	a_9)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_addr_0;
input 	a_9;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_13 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(a_9),
	.datab(seq_ac_addr_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'h5533;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_13 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_12 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_12 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_13 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_ba_0,
	ba_0)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_ba_0;
input 	ba_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x~1_combout ;
wire \ac_2x_2r~q ;
wire \ac_1t~q ;


altera_ddr_altddio_out_14 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(\ac_1t~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_add_1t_ac_lat_internal),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(seq_ac_ba_0),
	.datab(ba_0),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAACC;
defparam \ac_2x~1 .sum_lutc_input = "datac";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

endmodule

module altera_ddr_altddio_out_14 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_1jd auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_1jd (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_14 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_ba_1,
	ba_1)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_ba_1;
input 	ba_1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x~1_combout ;
wire \ac_2x_2r~q ;
wire \ac_1t~q ;


altera_ddr_altddio_out_15 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(\ac_1t~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_add_1t_ac_lat_internal),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(seq_ac_ba_1),
	.datab(ba_1),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAACC;
defparam \ac_2x~1 .sum_lutc_input = "datac";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

endmodule

module altera_ddr_altddio_out_15 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_1jd_1 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_1jd_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_15 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_cas_n_0,
	cas_n)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_cas_n_0;
input 	cas_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_16 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(gnd),
	.datab(ctl_init_success),
	.datac(seq_ac_cas_n_0),
	.datad(cas_n),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'hF3C0;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_16 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_13 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_13 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_16 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	ams_pipe_1,
	seq_ac_cke_0)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	ams_pipe_1;
input 	seq_ac_cke_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;
wire \ac_l~0_combout ;


altera_ddr_altddio_out_17 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.aclr(ams_pipe_1),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_1t~q ),
	.datab(ctl_init_success),
	.datac(seq_ac_cke_0),
	.datad(seq_ac_add_1t_ac_lat_internal),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hFAFC;
defparam \ac_2x~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(ctl_init_success),
	.datab(seq_ac_cke_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'hEEEE;
defparam \ac_l~0 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_17 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_1jd_2 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.aclr(aclr),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_1jd_2 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_17 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	ams_pipe_1,
	seq_ac_cs_n_0,
	cs_n_0)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	ams_pipe_1;
input 	seq_ac_cs_n_0;
input 	cs_n_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_18 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }),
	.aset(ams_pipe_1));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(gnd),
	.datab(ctl_init_success),
	.datac(seq_ac_cs_n_0),
	.datad(cs_n_0),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'hF3C0;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_18 (
	outclock,
	dataout,
	datain_l,
	datain_h,
	aset)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;
input 	aset;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_14 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}),
	.aset(aset));

endmodule

module altera_ddr_ddio_out_egd_14 (
	outclock,
	dataout,
	datain_l,
	datain_h,
	aset)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;
input 	aset;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(!aset),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_18 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_ras_n_0,
	ras_n)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_ras_n_0;
input 	ras_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_19 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(gnd),
	.datab(ctl_init_success),
	.datac(seq_ac_ras_n_0),
	.datad(ras_n),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'hF3C0;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_19 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_15 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_15 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ac_19 (
	phy_clk_1x,
	clk_2,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	seq_ac_we_n_0,
	we_n)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	clk_2;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	ctl_init_success;
input 	seq_ac_we_n_0;
input 	we_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_2x~q ;
wire \ac_2x_2r~q ;
wire \ac_l~0_combout ;
wire \ac_1t~q ;
wire \ac_2x~1_combout ;


altera_ddr_altddio_out_20 \full_rate.addr_pin (
	.outclock(clk_2),
	.dataout({dataout_0}),
	.datain_l({\ac_2x~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x(
	.clk(phy_clk_1x),
	.d(\ac_2x~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x~q ),
	.prn(vcc));
defparam ac_2x.is_wysiwyg = "true";
defparam ac_2x.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_2),
	.d(\ac_2x~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

cycloneiii_lcell_comb \ac_l~0 (
	.dataa(gnd),
	.datab(ctl_init_success),
	.datac(seq_ac_we_n_0),
	.datad(we_n),
	.cin(gnd),
	.combout(\ac_l~0_combout ),
	.cout());
defparam \ac_l~0 .lut_mask = 16'hF3C0;
defparam \ac_l~0 .sum_lutc_input = "datac";

dffeas ac_1t(
	.clk(phy_clk_1x),
	.d(\ac_l~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

cycloneiii_lcell_comb \ac_2x~1 (
	.dataa(\ac_l~0_combout ),
	.datab(gnd),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\ac_1t~q ),
	.cin(gnd),
	.combout(\ac_2x~1_combout ),
	.cout());
defparam \ac_2x~1 .lut_mask = 16'hAFA0;
defparam \ac_2x~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_out_20 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_out_egd_16 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module altera_ddr_ddio_out_egd_16 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_clk_reset (
	clk_0,
	clk_1,
	clk_2,
	clk_3,
	clk_4,
	ddio_outa_0,
	ddio_outa_01,
	reset_request_n,
	reset_phy_clk_1x_n1,
	ams_pipe_1,
	ams_pipe_11,
	seq_pll_inc_dec_n,
	seq_pll_start_reconfig,
	seq_mem_clk_disable,
	seq_pll_select,
	phs_shft_busy1,
	ams_pipe_12,
	input_cell_h_0,
	mem_clk_0,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=1 */;
output 	clk_0;
output 	clk_1;
output 	clk_2;
output 	clk_3;
output 	clk_4;
output 	ddio_outa_0;
output 	ddio_outa_01;
output 	reset_request_n;
output 	reset_phy_clk_1x_n1;
output 	ams_pipe_1;
output 	ams_pipe_11;
input 	seq_pll_inc_dec_n;
input 	seq_pll_start_reconfig;
input 	seq_mem_clk_disable;
input 	[2:0] seq_pll_select;
output 	phs_shft_busy1;
output 	ams_pipe_12;
output 	input_cell_h_0;
input 	mem_clk_0;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \pll|altpll_component|auto_generated|phasedone ;
wire \pll|altpll_component|auto_generated|pll1~LOCKED ;
wire \pll|altpll_component|auto_generated|pll_lock_sync~q ;
wire \pll_new_dir~q ;
wire \seq_pll_inc_dec_ccd~q ;
wire \pll_reprogram_request_pulse_2r~q ;
wire \pll_new_phase[0]~q ;
wire \pll_new_phase[1]~q ;
wire \pll_new_phase[2]~q ;
wire \always3~0_combout ;
wire \seq_pll_select_ccd[2]~q ;
wire \seq_pll_select_ccd[0]~q ;
wire \seq_pll_select_ccd[1]~q ;
wire \WideOr0~0_combout ;
wire \lookup~1_combout ;
wire \Decoder0~0_combout ;
wire \seq_pll_select_ccd[1]~0_combout ;
wire \phy_internal_reset_n~combout ;
wire \reset_master_ams~q ;
wire \global_pre_clear~q ;
wire \divider~5_combout ;
wire \phy_internal_reset_n~0_combout ;
wire \clk_div_reset_ams_n~q ;
wire \clk_div_reset_ams_n_r~q ;
wire \divider[0]~q ;
wire \divider[1]~4_combout ;
wire \divider[1]~q ;
wire \divider[2]~3_combout ;
wire \divider[2]~q ;
wire \scan_clk~2_combout ;
wire \scan_clk~q ;
wire \seq_pll_start_reconfig_ccd_pipe[0]~q ;
wire \seq_pll_start_reconfig_ccd_pipe[1]~q ;
wire \seq_pll_start_reconfig_ccd_pipe[2]~q ;
wire \pll_reconfig_reset_ams_n~q ;
wire \pll_reconfig_reset_ams_n_r~q ;
wire \seq_pll_start_reconfig_ams~q ;
wire \seq_pll_start_reconfig_r~q ;
wire \seq_pll_start_reconfig_2r~q ;
wire \seq_pll_start_reconfig_3r~q ;
wire \pll_phase_auto_calibrate_pulse~combout ;
wire \pll_reprogram_request_pulse~q ;
wire \pll_reprogram_request_pulse_r~q ;
wire \pll_reprogram_request_long_pulse~1_combout ;
wire \pll_reprogram_request~q ;
wire \phs_shft_busy~0_combout ;


altera_ddr_altera_ddr_phy_alt_mem_phy_pll pll(
	.phasedone(\pll|altpll_component|auto_generated|phasedone ),
	.pll1(\pll|altpll_component|auto_generated|pll1~LOCKED ),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_2(clk_2),
	.clk_3(clk_3),
	.clk_4(clk_4),
	.pll_lock_sync(\pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.locked(reset_request_n),
	.pll_new_dir(\pll_new_dir~q ),
	.pll_reprogram_request(\pll_reprogram_request~q ),
	.scan_clk(\scan_clk~q ),
	.pll_new_phase_0(\pll_new_phase[0]~q ),
	.pll_new_phase_1(\pll_new_phase[1]~q ),
	.pll_new_phase_2(\pll_new_phase[2]~q ),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk));

altera_ddr_altddio_bidir_2 \DDR_CLK_OUT[0].ddr_clk_out_p (
	.outclock(clk_1),
	.inclock(clk_4),
	.ddio_outa_0(ddio_outa_0),
	.aclr(seq_mem_clk_disable),
	.input_cell_h_0(input_cell_h_0),
	.mem_clk_0(mem_clk_0));

altera_ddr_altddio_bidir_1 \DDR_CLK_OUT[0].ddr_clk_out_n (
	.outclock(clk_1),
	.ddio_outa_0(ddio_outa_01),
	.aclr(seq_mem_clk_disable));

altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe ac_clk_pipe_2x(
	.clock(clk_2),
	.ams_pipe_1(ams_pipe_1),
	.pre_clear(\global_pre_clear~q ));

altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe_2 measure_clk_pipe(
	.clock(clk_4),
	.pre_clear(\global_pre_clear~q ),
	.ams_pipe_1(ams_pipe_12));

altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe_6 resync_clk_pipe(
	.clock(clk_3),
	.pre_clear(\global_pre_clear~q ),
	.ams_pipe_1(ams_pipe_11));

dffeas pll_new_dir(
	.clk(\scan_clk~q ),
	.d(\seq_pll_inc_dec_ccd~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_dir~q ),
	.prn(vcc));
defparam pll_new_dir.is_wysiwyg = "true";
defparam pll_new_dir.power_up = "low";

dffeas seq_pll_inc_dec_ccd(
	.clk(clk_1),
	.d(seq_pll_inc_dec_n),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_inc_dec_ccd~q ),
	.prn(vcc));
defparam seq_pll_inc_dec_ccd.is_wysiwyg = "true";
defparam seq_pll_inc_dec_ccd.power_up = "low";

dffeas pll_reprogram_request_pulse_2r(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_pulse_r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse_2r~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse_2r.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse_2r.power_up = "low";

dffeas \pll_new_phase[0] (
	.clk(\scan_clk~q ),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[0]~q ),
	.prn(vcc));
defparam \pll_new_phase[0] .is_wysiwyg = "true";
defparam \pll_new_phase[0] .power_up = "low";

dffeas \pll_new_phase[1] (
	.clk(\scan_clk~q ),
	.d(\lookup~1_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[1]~q ),
	.prn(vcc));
defparam \pll_new_phase[1] .is_wysiwyg = "true";
defparam \pll_new_phase[1] .power_up = "low";

dffeas \pll_new_phase[2] (
	.clk(\scan_clk~q ),
	.d(\Decoder0~0_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[2]~q ),
	.prn(vcc));
defparam \pll_new_phase[2] .is_wysiwyg = "true";
defparam \pll_new_phase[2] .power_up = "low";

cycloneiii_lcell_comb \always3~0 (
	.dataa(seq_pll_start_reconfig),
	.datab(gnd),
	.datac(gnd),
	.datad(\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hAAFF;
defparam \always3~0 .sum_lutc_input = "datac";

dffeas \seq_pll_select_ccd[2] (
	.clk(clk_1),
	.d(seq_pll_select[2]),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[2]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[2] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[2] .power_up = "low";

dffeas \seq_pll_select_ccd[0] (
	.clk(clk_1),
	.d(seq_pll_select[0]),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[0]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[0] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[0] .power_up = "low";

dffeas \seq_pll_select_ccd[1] (
	.clk(clk_1),
	.d(\seq_pll_select_ccd[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[1]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[1] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[1] .power_up = "low";

cycloneiii_lcell_comb \WideOr0~0 (
	.dataa(\seq_pll_select_ccd[2]~q ),
	.datab(gnd),
	.datac(\seq_pll_select_ccd[0]~q ),
	.datad(\seq_pll_select_ccd[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hAFFA;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \lookup~1 (
	.dataa(\seq_pll_select_ccd[1]~q ),
	.datab(\seq_pll_select_ccd[2]~q ),
	.datac(gnd),
	.datad(\seq_pll_select_ccd[0]~q ),
	.cin(gnd),
	.combout(\lookup~1_combout ),
	.cout());
defparam \lookup~1 .lut_mask = 16'h66FF;
defparam \lookup~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Decoder0~0 (
	.dataa(\seq_pll_select_ccd[1]~q ),
	.datab(\seq_pll_select_ccd[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
defparam \Decoder0~0 .lut_mask = 16'hEEEE;
defparam \Decoder0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_select_ccd[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_pll_select_ccd[1]~0_combout ),
	.cout());
defparam \seq_pll_select_ccd[1]~0 .lut_mask = 16'h0000;
defparam \seq_pll_select_ccd[1]~0 .sum_lutc_input = "datac";

dffeas reset_phy_clk_1x_n(
	.clk(clk_1),
	.d(vcc),
	.asdata(vcc),
	.clrn(\global_pre_clear~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_phy_clk_1x_n1),
	.prn(vcc));
defparam reset_phy_clk_1x_n.is_wysiwyg = "true";
defparam reset_phy_clk_1x_n.power_up = "low";

dffeas phs_shft_busy(
	.clk(\scan_clk~q ),
	.d(\phs_shft_busy~0_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(phs_shft_busy1),
	.prn(vcc));
defparam phs_shft_busy.is_wysiwyg = "true";
defparam phs_shft_busy.power_up = "low";

cycloneiii_lcell_comb phy_internal_reset_n(
	.dataa(\pll|altpll_component|auto_generated|pll1~LOCKED ),
	.datab(\pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.datac(global_reset_n),
	.datad(soft_reset_n),
	.cin(gnd),
	.combout(\phy_internal_reset_n~combout ),
	.cout());
defparam phy_internal_reset_n.lut_mask = 16'h7FFF;
defparam phy_internal_reset_n.sum_lutc_input = "datac";

dffeas reset_master_ams(
	.clk(clk_1),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_master_ams~q ),
	.prn(vcc));
defparam reset_master_ams.is_wysiwyg = "true";
defparam reset_master_ams.power_up = "low";

dffeas global_pre_clear(
	.clk(clk_1),
	.d(\reset_master_ams~q ),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\global_pre_clear~q ),
	.prn(vcc));
defparam global_pre_clear.is_wysiwyg = "true";
defparam global_pre_clear.power_up = "low";

cycloneiii_lcell_comb \divider~5 (
	.dataa(\divider[0]~q ),
	.datab(gnd),
	.datac(\divider[2]~q ),
	.datad(\divider[1]~q ),
	.cin(gnd),
	.combout(\divider~5_combout ),
	.cout());
defparam \divider~5 .lut_mask = 16'hFFF5;
defparam \divider~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \phy_internal_reset_n~0 (
	.dataa(\pll|altpll_component|auto_generated|pll1~LOCKED ),
	.datab(\pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.datac(global_reset_n),
	.datad(gnd),
	.cin(gnd),
	.combout(\phy_internal_reset_n~0_combout ),
	.cout());
defparam \phy_internal_reset_n~0 .lut_mask = 16'h7F7F;
defparam \phy_internal_reset_n~0 .sum_lutc_input = "datac";

dffeas clk_div_reset_ams_n(
	.clk(clk_1),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_div_reset_ams_n~q ),
	.prn(vcc));
defparam clk_div_reset_ams_n.is_wysiwyg = "true";
defparam clk_div_reset_ams_n.power_up = "low";

dffeas clk_div_reset_ams_n_r(
	.clk(clk_1),
	.d(\clk_div_reset_ams_n~q ),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_div_reset_ams_n_r~q ),
	.prn(vcc));
defparam clk_div_reset_ams_n_r.is_wysiwyg = "true";
defparam clk_div_reset_ams_n_r.power_up = "low";

dffeas \divider[0] (
	.clk(clk_1),
	.d(\divider~5_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[0]~q ),
	.prn(vcc));
defparam \divider[0] .is_wysiwyg = "true";
defparam \divider[0] .power_up = "low";

cycloneiii_lcell_comb \divider[1]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\divider[1]~q ),
	.datad(\divider[0]~q ),
	.cin(gnd),
	.combout(\divider[1]~4_combout ),
	.cout());
defparam \divider[1]~4 .lut_mask = 16'h0FF0;
defparam \divider[1]~4 .sum_lutc_input = "datac";

dffeas \divider[1] (
	.clk(clk_1),
	.d(\divider[1]~4_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[1]~q ),
	.prn(vcc));
defparam \divider[1] .is_wysiwyg = "true";
defparam \divider[1] .power_up = "low";

cycloneiii_lcell_comb \divider[2]~3 (
	.dataa(gnd),
	.datab(\divider[2]~q ),
	.datac(\divider[1]~q ),
	.datad(\divider[0]~q ),
	.cin(gnd),
	.combout(\divider[2]~3_combout ),
	.cout());
defparam \divider[2]~3 .lut_mask = 16'hC33C;
defparam \divider[2]~3 .sum_lutc_input = "datac";

dffeas \divider[2] (
	.clk(clk_1),
	.d(\divider[2]~3_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[2]~q ),
	.prn(vcc));
defparam \divider[2] .is_wysiwyg = "true";
defparam \divider[2] .power_up = "low";

cycloneiii_lcell_comb \scan_clk~2 (
	.dataa(\scan_clk~q ),
	.datab(\divider[2]~q ),
	.datac(\divider[1]~q ),
	.datad(\divider[0]~q ),
	.cin(gnd),
	.combout(\scan_clk~2_combout ),
	.cout());
defparam \scan_clk~2 .lut_mask = 16'h6996;
defparam \scan_clk~2 .sum_lutc_input = "datac";

dffeas scan_clk(
	.clk(clk_1),
	.d(\scan_clk~2_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_clk~q ),
	.prn(vcc));
defparam scan_clk.is_wysiwyg = "true";
defparam scan_clk.power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[0] (
	.clk(clk_1),
	.d(seq_pll_start_reconfig),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[0] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[0] .power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[1] (
	.clk(clk_1),
	.d(\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[1]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[1] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[1] .power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[2] (
	.clk(clk_1),
	.d(\seq_pll_start_reconfig_ccd_pipe[1]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[2]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[2] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[2] .power_up = "low";

dffeas pll_reconfig_reset_ams_n(
	.clk(\scan_clk~q ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reconfig_reset_ams_n~q ),
	.prn(vcc));
defparam pll_reconfig_reset_ams_n.is_wysiwyg = "true";
defparam pll_reconfig_reset_ams_n.power_up = "low";

dffeas pll_reconfig_reset_ams_n_r(
	.clk(\scan_clk~q ),
	.d(\pll_reconfig_reset_ams_n~q ),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reconfig_reset_ams_n_r~q ),
	.prn(vcc));
defparam pll_reconfig_reset_ams_n_r.is_wysiwyg = "true";
defparam pll_reconfig_reset_ams_n_r.power_up = "low";

dffeas seq_pll_start_reconfig_ams(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_ccd_pipe[2]~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ams~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_ams.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_ams.power_up = "low";

dffeas seq_pll_start_reconfig_r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_ams~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_r.power_up = "low";

dffeas seq_pll_start_reconfig_2r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_2r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_2r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_2r.power_up = "low";

dffeas seq_pll_start_reconfig_3r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_2r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_3r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_3r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_3r.power_up = "low";

cycloneiii_lcell_comb pll_phase_auto_calibrate_pulse(
	.dataa(\seq_pll_start_reconfig_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\seq_pll_start_reconfig_3r~q ),
	.cin(gnd),
	.combout(\pll_phase_auto_calibrate_pulse~combout ),
	.cout());
defparam pll_phase_auto_calibrate_pulse.lut_mask = 16'hAAFF;
defparam pll_phase_auto_calibrate_pulse.sum_lutc_input = "datac";

dffeas pll_reprogram_request_pulse(
	.clk(\scan_clk~q ),
	.d(\pll_phase_auto_calibrate_pulse~combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse.power_up = "low";

dffeas pll_reprogram_request_pulse_r(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_pulse~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse_r~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse_r.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse_r.power_up = "low";

cycloneiii_lcell_comb \pll_reprogram_request_long_pulse~1 (
	.dataa(\pll_reprogram_request_pulse_2r~q ),
	.datab(\pll_reprogram_request_pulse~q ),
	.datac(\pll_reprogram_request_pulse_r~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pll_reprogram_request_long_pulse~1_combout ),
	.cout());
defparam \pll_reprogram_request_long_pulse~1 .lut_mask = 16'hFEFE;
defparam \pll_reprogram_request_long_pulse~1 .sum_lutc_input = "datac";

dffeas pll_reprogram_request(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_long_pulse~1_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request~q ),
	.prn(vcc));
defparam pll_reprogram_request.is_wysiwyg = "true";
defparam pll_reprogram_request.power_up = "low";

cycloneiii_lcell_comb \phs_shft_busy~0 (
	.dataa(\pll_reprogram_request~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\pll|altpll_component|auto_generated|phasedone ),
	.cin(gnd),
	.combout(\phs_shft_busy~0_combout ),
	.cout());
defparam \phs_shft_busy~0 .lut_mask = 16'hAAFF;
defparam \phs_shft_busy~0 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altddio_bidir_1 (
	outclock,
	ddio_outa_0,
	aclr)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	ddio_outa_0;
input 	aclr;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_bidir_idf auto_generated(
	.outclock(outclock),
	.ddio_outa_0(ddio_outa_0),
	.aclr(aclr));

endmodule

module altera_ddr_ddio_bidir_idf (
	outclock,
	ddio_outa_0,
	aclr)/* synthesis synthesis_greybox=1 */;
input 	outclock;
output 	ddio_outa_0;
input 	aclr;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(vcc),
	.datainhi(gnd),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.dataout(ddio_outa_0),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module altera_ddr_altddio_bidir_2 (
	outclock,
	inclock,
	ddio_outa_0,
	aclr,
	input_cell_h_0,
	mem_clk_0)/* synthesis synthesis_greybox=1 */;
input 	outclock;
input 	inclock;
output 	ddio_outa_0;
input 	aclr;
output 	input_cell_h_0;
input 	mem_clk_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_bidir_e4h auto_generated(
	.outclock(outclock),
	.inclock(inclock),
	.ddio_outa_0(ddio_outa_0),
	.aclr(aclr),
	.input_cell_h_0(input_cell_h_0),
	.mem_clk_0(mem_clk_0));

endmodule

module altera_ddr_ddio_bidir_e4h (
	outclock,
	inclock,
	ddio_outa_0,
	aclr,
	input_cell_h_0,
	mem_clk_0)/* synthesis synthesis_greybox=1 */;
input 	outclock;
input 	inclock;
output 	ddio_outa_0;
input 	aclr;
output 	input_cell_h_0;
input 	mem_clk_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_ddio_out \ddio_outa[0] (
	.datainlo(vcc),
	.datainhi(gnd),
	.clkhi(!outclock),
	.clklo(!outclock),
	.muxsel(!outclock),
	.clk(gnd),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.dataout(ddio_outa_0),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(mem_clk_0),
	.asdata(vcc),
	.clrn(aclr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_pll (
	phasedone,
	pll1,
	clk_0,
	clk_1,
	clk_2,
	clk_3,
	clk_4,
	pll_lock_sync,
	locked,
	pll_new_dir,
	pll_reprogram_request,
	scan_clk,
	pll_new_phase_0,
	pll_new_phase_1,
	pll_new_phase_2,
	global_reset_n,
	pll_ref_clk)/* synthesis synthesis_greybox=1 */;
output 	phasedone;
output 	pll1;
output 	clk_0;
output 	clk_1;
output 	clk_2;
output 	clk_3;
output 	clk_4;
output 	pll_lock_sync;
output 	locked;
input 	pll_new_dir;
input 	pll_reprogram_request;
input 	scan_clk;
input 	pll_new_phase_0;
input 	pll_new_phase_1;
input 	pll_new_phase_2;
input 	global_reset_n;
input 	pll_ref_clk;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altpll_1 altpll_component(
	.phasedone(phasedone),
	.pll1(pll1),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_2(clk_2),
	.clk_3(clk_3),
	.clk_4(clk_4),
	.pll_lock_sync(pll_lock_sync),
	.locked(locked),
	.phaseupdown(pll_new_dir),
	.phasestep(pll_reprogram_request),
	.scanclk(scan_clk),
	.pll_new_phase_0(pll_new_phase_0),
	.pll_new_phase_1(pll_new_phase_1),
	.pll_new_phase_2(pll_new_phase_2),
	.areset(global_reset_n),
	.inclk({gnd,pll_ref_clk}));

endmodule

module altera_ddr_altpll_1 (
	phasedone,
	pll1,
	clk_0,
	clk_1,
	clk_2,
	clk_3,
	clk_4,
	pll_lock_sync,
	locked,
	phaseupdown,
	phasestep,
	scanclk,
	pll_new_phase_0,
	pll_new_phase_1,
	pll_new_phase_2,
	areset,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	phasedone;
output 	pll1;
output 	clk_0;
output 	clk_1;
output 	clk_2;
output 	clk_3;
output 	clk_4;
output 	pll_lock_sync;
output 	locked;
input 	phaseupdown;
input 	phasestep;
input 	scanclk;
input 	pll_new_phase_0;
input 	pll_new_phase_1;
input 	pll_new_phase_2;
input 	areset;
input 	[1:0] inclk;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altpll_8g53 auto_generated(
	.phasedone(phasedone),
	.pll11(pll1),
	.clk({clk_4,clk_3,clk_2,clk_1,clk_0}),
	.pll_lock_sync1(pll_lock_sync),
	.locked1(locked),
	.phaseupdown(phaseupdown),
	.phasestep(phasestep),
	.scanclk(scanclk),
	.pll_new_phase_0(pll_new_phase_0),
	.pll_new_phase_1(pll_new_phase_1),
	.pll_new_phase_2(pll_new_phase_2),
	.areset(areset),
	.inclk({gnd,inclk[0]}));

endmodule

module altera_ddr_altpll_8g53 (
	phasedone,
	pll11,
	clk,
	pll_lock_sync1,
	locked1,
	phaseupdown,
	phasestep,
	scanclk,
	pll_new_phase_0,
	pll_new_phase_1,
	pll_new_phase_2,
	areset,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	phasedone;
output 	pll11;
output 	[4:0] clk;
output 	pll_lock_sync1;
output 	locked1;
input 	phaseupdown;
input 	phasestep;
input 	scanclk;
input 	pll_new_phase_0;
input 	pll_new_phase_1;
input 	pll_new_phase_2;
input 	areset;
input 	[1:0] inclk;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \altpll_dyn_phase_le2|combout ;
wire \altpll_dyn_phase_le4|combout ;
wire \altpll_dyn_phase_le5|combout ;
wire \remap_decoy_le3a[0]~combout ;
wire \remap_decoy_le3a[1]~combout ;
wire \remap_decoy_le3a[2]~combout ;
wire \pll1~FBOUT ;

wire [4:0] pll1_CLK_bus;

assign clk[0] = pll1_CLK_bus[0];
assign clk[1] = pll1_CLK_bus[1];
assign clk[2] = pll1_CLK_bus[2];
assign clk[3] = pll1_CLK_bus[3];
assign clk[4] = pll1_CLK_bus[4];

altera_ddr_altpll_dyn_phase_le_9ii altpll_dyn_phase_le2(
	.combout(\altpll_dyn_phase_le2|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ));

altera_ddr_altpll_dyn_phase_le_aii altpll_dyn_phase_le4(
	.combout(\altpll_dyn_phase_le4|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ));

altera_ddr_altpll_dyn_phase_le_bii altpll_dyn_phase_le5(
	.combout(\altpll_dyn_phase_le5|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ));

cycloneiii_lcell_comb \remap_decoy_le3a[0] (
	.dataa(pll_new_phase_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\remap_decoy_le3a[0]~combout ),
	.cout());
defparam \remap_decoy_le3a[0] .lut_mask = 16'hAAAA;
defparam \remap_decoy_le3a[0] .sum_lutc_input = "datac";

cycloneiii_lcell_comb \remap_decoy_le3a[1] (
	.dataa(pll_new_phase_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\remap_decoy_le3a[1]~combout ),
	.cout());
defparam \remap_decoy_le3a[1] .lut_mask = 16'hAAAA;
defparam \remap_decoy_le3a[1] .sum_lutc_input = "datac";

cycloneiii_lcell_comb \remap_decoy_le3a[2] (
	.dataa(pll_new_phase_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\remap_decoy_le3a[2]~combout ),
	.cout());
defparam \remap_decoy_le3a[2] .lut_mask = 16'hAAAA;
defparam \remap_decoy_le3a[2] .sum_lutc_input = "datac";

cycloneiii_pll pll1(
	.areset(!areset),
	.pfdena(vcc),
	.fbin(\pll1~FBOUT ),
	.phaseupdown(phaseupdown),
	.phasestep(phasestep),
	.scandata(gnd),
	.scanclk(scanclk),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect({\altpll_dyn_phase_le5|combout ,\altpll_dyn_phase_le4|combout ,\altpll_dyn_phase_le2|combout }),
	.phasedone(phasedone),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(pll11),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(\pll1~FBOUT ),
	.clk(pll1_CLK_bus),
	.clkbad());
defparam pll1.auto_settings = "false";
defparam pll1.bandwidth_type = "auto";
defparam pll1.c0_high = 8;
defparam pll1.c0_initial = 3;
defparam pll1.c0_low = 8;
defparam pll1.c0_mode = "even";
defparam pll1.c0_ph = 0;
defparam pll1.c1_high = 4;
defparam pll1.c1_initial = 3;
defparam pll1.c1_low = 4;
defparam pll1.c1_mode = "even";
defparam pll1.c1_ph = 0;
defparam pll1.c1_use_casc_in = "off";
defparam pll1.c2_high = 4;
defparam pll1.c2_initial = 1;
defparam pll1.c2_low = 4;
defparam pll1.c2_mode = "even";
defparam pll1.c2_ph = 0;
defparam pll1.c2_use_casc_in = "off";
defparam pll1.c3_high = 4;
defparam pll1.c3_initial = 3;
defparam pll1.c3_low = 4;
defparam pll1.c3_mode = "even";
defparam pll1.c3_ph = 0;
defparam pll1.c3_use_casc_in = "off";
defparam pll1.c4_high = 4;
defparam pll1.c4_initial = 3;
defparam pll1.c4_low = 4;
defparam pll1.c4_mode = "even";
defparam pll1.c4_ph = 0;
defparam pll1.c4_use_casc_in = "off";
defparam pll1.charge_pump_current_bits = 1;
defparam pll1.clk0_counter = "c0";
defparam pll1.clk0_divide_by = 2;
defparam pll1.clk0_duty_cycle = 50;
defparam pll1.clk0_multiply_by = 3;
defparam pll1.clk0_phase_shift = "0";
defparam pll1.clk1_counter = "c1";
defparam pll1.clk1_divide_by = 1;
defparam pll1.clk1_duty_cycle = 50;
defparam pll1.clk1_multiply_by = 3;
defparam pll1.clk1_phase_shift = "0";
defparam pll1.clk2_counter = "c2";
defparam pll1.clk2_divide_by = 1;
defparam pll1.clk2_duty_cycle = 50;
defparam pll1.clk2_multiply_by = 3;
defparam pll1.clk2_phase_shift = "-1667";
defparam pll1.clk3_counter = "c3";
defparam pll1.clk3_divide_by = 1;
defparam pll1.clk3_duty_cycle = 50;
defparam pll1.clk3_multiply_by = 3;
defparam pll1.clk3_phase_shift = "0";
defparam pll1.clk4_counter = "c4";
defparam pll1.clk4_divide_by = 1;
defparam pll1.clk4_duty_cycle = 50;
defparam pll1.clk4_multiply_by = 3;
defparam pll1.clk4_phase_shift = "0";
defparam pll1.compensate_clock = "clock1";
defparam pll1.inclk0_input_frequency = 20000;
defparam pll1.inclk1_input_frequency = 0;
defparam pll1.loop_filter_c_bits = 0;
defparam pll1.loop_filter_r_bits = 27;
defparam pll1.m = 24;
defparam pll1.m_initial = 3;
defparam pll1.m_ph = 0;
defparam pll1.n = 1;
defparam pll1.operation_mode = "normal";
defparam pll1.pfd_max = 200000;
defparam pll1.pfd_min = 3076;
defparam pll1.self_reset_on_loss_lock = "off";
defparam pll1.simulation_type = "timing";
defparam pll1.switch_over_type = "auto";
defparam pll1.vco_center = 769;
defparam pll1.vco_divide_by = 0;
defparam pll1.vco_frequency_control = "auto";
defparam pll1.vco_max = 1666;
defparam pll1.vco_min = 769;
defparam pll1.vco_multiply_by = 0;
defparam pll1.vco_phase_shift_step = 104;
defparam pll1.vco_post_scale = 1;

dffeas pll_lock_sync(
	.clk(pll11),
	.d(vcc),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pll_lock_sync1),
	.prn(vcc));
defparam pll_lock_sync.is_wysiwyg = "true";
defparam pll_lock_sync.power_up = "low";

cycloneiii_lcell_comb locked(
	.dataa(pll11),
	.datab(pll_lock_sync1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(locked1),
	.cout());
defparam locked.lut_mask = 16'hEEEE;
defparam locked.sum_lutc_input = "datac";

endmodule

module altera_ddr_altpll_dyn_phase_le_9ii (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2)/* synthesis synthesis_greybox=1 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_lcell_comb le_comb6(
	.dataa(remap_decoy_le3a_0),
	.datab(remap_decoy_le3a_1),
	.datac(remap_decoy_le3a_2),
	.datad(gnd),
	.cin(gnd),
	.combout(combout),
	.cout());
defparam le_comb6.lut_mask = 16'hAAAA;
defparam le_comb6.sum_lutc_input = "datac";

endmodule

module altera_ddr_altpll_dyn_phase_le_aii (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2)/* synthesis synthesis_greybox=1 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_lcell_comb le_comb7(
	.dataa(remap_decoy_le3a_0),
	.datab(remap_decoy_le3a_1),
	.datac(remap_decoy_le3a_2),
	.datad(gnd),
	.cin(gnd),
	.combout(combout),
	.cout());
defparam le_comb7.lut_mask = 16'hCCCC;
defparam le_comb7.sum_lutc_input = "datac";

endmodule

module altera_ddr_altpll_dyn_phase_le_bii (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2)/* synthesis synthesis_greybox=1 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



cycloneiii_lcell_comb le_comb8(
	.dataa(remap_decoy_le3a_0),
	.datab(remap_decoy_le3a_1),
	.datac(remap_decoy_le3a_2),
	.datad(gnd),
	.cin(gnd),
	.combout(combout),
	.cout());
defparam le_comb8.lut_mask = 16'hF0F0;
defparam le_comb8.sum_lutc_input = "datac";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe (
	clock,
	ams_pipe_1,
	pre_clear)/* synthesis synthesis_greybox=1 */;
input 	clock;
output 	ams_pipe_1;
input 	pre_clear;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe_2 (
	clock,
	pre_clear,
	ams_pipe_1)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	pre_clear;
output 	ams_pipe_1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_reset_pipe_6 (
	clock,
	pre_clear,
	ams_pipe_1)/* synthesis synthesis_greybox=1 */;
input 	clock;
input 	pre_clear;
output 	ams_pipe_1;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_dp_io (
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	mem_clk_2x,
	write_clk_2x,
	clk_3,
	dm_ddio_dataout_0,
	dm_ddio_dataout_1,
	dq_ddio_dataout_0,
	dq_ddio_dataout_1,
	dq_ddio_dataout_2,
	dq_ddio_dataout_3,
	dq_ddio_dataout_4,
	dq_ddio_dataout_5,
	dq_ddio_dataout_6,
	dq_ddio_dataout_7,
	dq_ddio_dataout_8,
	dq_ddio_dataout_9,
	dq_ddio_dataout_10,
	dq_ddio_dataout_11,
	dq_ddio_dataout_12,
	dq_ddio_dataout_13,
	dq_ddio_dataout_14,
	dq_ddio_dataout_15,
	dqs_ddio_dataout_0,
	wdp_wdqs_oe_2x_r_0,
	dqs_ddio_dataout_1,
	wdp_wdqs_oe_2x_r_1,
	wdp_dm_l_2x,
	wdp_dm_h_2x,
	ams_pipe_1,
	wdp_wdata_oe_2x_r_0,
	wdp_wdata_oe_2x_r_1,
	wdp_wdata_oe_2x_r_2,
	wdp_wdata_oe_2x_r_3,
	wdp_wdata_oe_2x_r_4,
	wdp_wdata_oe_2x_r_5,
	wdp_wdata_oe_2x_r_6,
	wdp_wdata_oe_2x_r_7,
	wdp_wdata_oe_2x_r_8,
	wdp_wdata_oe_2x_r_9,
	wdp_wdata_oe_2x_r_10,
	wdp_wdata_oe_2x_r_11,
	wdp_wdata_oe_2x_r_12,
	wdp_wdata_oe_2x_r_13,
	wdp_wdata_oe_2x_r_14,
	wdp_wdata_oe_2x_r_15,
	dio_rdata_h_2x_0,
	dio_rdata_h_2x_1,
	dio_rdata_h_2x_2,
	dio_rdata_h_2x_3,
	dio_rdata_h_2x_4,
	dio_rdata_h_2x_5,
	dio_rdata_h_2x_6,
	dio_rdata_h_2x_7,
	dio_rdata_h_2x_8,
	dio_rdata_h_2x_9,
	dio_rdata_h_2x_10,
	dio_rdata_h_2x_11,
	dio_rdata_h_2x_12,
	dio_rdata_h_2x_13,
	dio_rdata_h_2x_14,
	dio_rdata_h_2x_15,
	dio_rdata_l_2x_0,
	dio_rdata_l_2x_1,
	dio_rdata_l_2x_2,
	dio_rdata_l_2x_3,
	dio_rdata_l_2x_4,
	dio_rdata_l_2x_5,
	dio_rdata_l_2x_6,
	dio_rdata_l_2x_7,
	dio_rdata_l_2x_8,
	dio_rdata_l_2x_9,
	dio_rdata_l_2x_10,
	dio_rdata_l_2x_11,
	dio_rdata_l_2x_12,
	dio_rdata_l_2x_13,
	dio_rdata_l_2x_14,
	dio_rdata_l_2x_15,
	wdp_wdata_l_2x,
	wdp_wdata_h_2x,
	wdp_wdata_oe_2x,
	wdp_wdqs_2x,
	wdp_wdqs_oe_2x)/* synthesis synthesis_greybox=1 */;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
input 	mem_clk_2x;
input 	write_clk_2x;
input 	clk_3;
output 	dm_ddio_dataout_0;
output 	dm_ddio_dataout_1;
output 	dq_ddio_dataout_0;
output 	dq_ddio_dataout_1;
output 	dq_ddio_dataout_2;
output 	dq_ddio_dataout_3;
output 	dq_ddio_dataout_4;
output 	dq_ddio_dataout_5;
output 	dq_ddio_dataout_6;
output 	dq_ddio_dataout_7;
output 	dq_ddio_dataout_8;
output 	dq_ddio_dataout_9;
output 	dq_ddio_dataout_10;
output 	dq_ddio_dataout_11;
output 	dq_ddio_dataout_12;
output 	dq_ddio_dataout_13;
output 	dq_ddio_dataout_14;
output 	dq_ddio_dataout_15;
output 	dqs_ddio_dataout_0;
output 	wdp_wdqs_oe_2x_r_0;
output 	dqs_ddio_dataout_1;
output 	wdp_wdqs_oe_2x_r_1;
input 	[1:0] wdp_dm_l_2x;
input 	[1:0] wdp_dm_h_2x;
input 	ams_pipe_1;
output 	wdp_wdata_oe_2x_r_0;
output 	wdp_wdata_oe_2x_r_1;
output 	wdp_wdata_oe_2x_r_2;
output 	wdp_wdata_oe_2x_r_3;
output 	wdp_wdata_oe_2x_r_4;
output 	wdp_wdata_oe_2x_r_5;
output 	wdp_wdata_oe_2x_r_6;
output 	wdp_wdata_oe_2x_r_7;
output 	wdp_wdata_oe_2x_r_8;
output 	wdp_wdata_oe_2x_r_9;
output 	wdp_wdata_oe_2x_r_10;
output 	wdp_wdata_oe_2x_r_11;
output 	wdp_wdata_oe_2x_r_12;
output 	wdp_wdata_oe_2x_r_13;
output 	wdp_wdata_oe_2x_r_14;
output 	wdp_wdata_oe_2x_r_15;
output 	dio_rdata_h_2x_0;
output 	dio_rdata_h_2x_1;
output 	dio_rdata_h_2x_2;
output 	dio_rdata_h_2x_3;
output 	dio_rdata_h_2x_4;
output 	dio_rdata_h_2x_5;
output 	dio_rdata_h_2x_6;
output 	dio_rdata_h_2x_7;
output 	dio_rdata_h_2x_8;
output 	dio_rdata_h_2x_9;
output 	dio_rdata_h_2x_10;
output 	dio_rdata_h_2x_11;
output 	dio_rdata_h_2x_12;
output 	dio_rdata_h_2x_13;
output 	dio_rdata_h_2x_14;
output 	dio_rdata_h_2x_15;
output 	dio_rdata_l_2x_0;
output 	dio_rdata_l_2x_1;
output 	dio_rdata_l_2x_2;
output 	dio_rdata_l_2x_3;
output 	dio_rdata_l_2x_4;
output 	dio_rdata_l_2x_5;
output 	dio_rdata_l_2x_6;
output 	dio_rdata_l_2x_7;
output 	dio_rdata_l_2x_8;
output 	dio_rdata_l_2x_9;
output 	dio_rdata_l_2x_10;
output 	dio_rdata_l_2x_11;
output 	dio_rdata_l_2x_12;
output 	dio_rdata_l_2x_13;
output 	dio_rdata_l_2x_14;
output 	dio_rdata_l_2x_15;
input 	[15:0] wdp_wdata_l_2x;
input 	[15:0] wdp_wdata_h_2x;
input 	[15:0] wdp_wdata_oe_2x;
input 	[1:0] wdp_wdqs_2x;
input 	[1:0] wdp_wdqs_oe_2x;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \dqs_group[0].dq[0].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[1].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[2].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[3].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[4].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[5].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[6].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[7].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[0].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[1].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[2].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[3].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[4].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[5].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[6].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[1].dq[7].dqi|auto_generated|input_latch_l[0]~q ;
wire \dqs_group[0].dq[0].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[1].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[2].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[3].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[4].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[5].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[6].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[0].dq[7].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[0].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[1].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[2].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[3].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[4].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[5].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[6].dqi|auto_generated|input_cell_h[0]~q ;
wire \dqs_group[1].dq[7].dqi|auto_generated|input_cell_h[0]~q ;
wire \rdata_p_ams[0]~q ;
wire \rdata_p_ams[1]~q ;
wire \rdata_p_ams[2]~q ;
wire \rdata_p_ams[3]~q ;
wire \rdata_p_ams[4]~q ;
wire \rdata_p_ams[5]~q ;
wire \rdata_p_ams[6]~q ;
wire \rdata_p_ams[7]~q ;
wire \rdata_p_ams[8]~q ;
wire \rdata_p_ams[9]~q ;
wire \rdata_p_ams[10]~q ;
wire \rdata_p_ams[11]~q ;
wire \rdata_p_ams[12]~q ;
wire \rdata_p_ams[13]~q ;
wire \rdata_p_ams[14]~q ;
wire \rdata_p_ams[15]~q ;
wire \rdata_n_ams[0]~q ;
wire \rdata_n_ams[1]~q ;
wire \rdata_n_ams[2]~q ;
wire \rdata_n_ams[3]~q ;
wire \rdata_n_ams[4]~q ;
wire \rdata_n_ams[5]~q ;
wire \rdata_n_ams[6]~q ;
wire \rdata_n_ams[7]~q ;
wire \rdata_n_ams[8]~q ;
wire \rdata_n_ams[9]~q ;
wire \rdata_n_ams[10]~q ;
wire \rdata_n_ams[11]~q ;
wire \rdata_n_ams[12]~q ;
wire \rdata_n_ams[13]~q ;
wire \rdata_n_ams[14]~q ;
wire \rdata_n_ams[15]~q ;


altera_ddr_altddio_in_1 \dqs_group[0].dq[0].dqi (
	.datain({dq_datain_0}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[0].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[0].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_2 \dqs_group[0].dq[1].dqi (
	.datain({dq_datain_1}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[1].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[1].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_3 \dqs_group[0].dq[2].dqi (
	.datain({dq_datain_2}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[2].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[2].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_4 \dqs_group[0].dq[3].dqi (
	.datain({dq_datain_3}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[3].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[3].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_5 \dqs_group[0].dq[4].dqi (
	.datain({dq_datain_4}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[4].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[4].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_6 \dqs_group[0].dq[5].dqi (
	.datain({dq_datain_5}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[5].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[5].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_7 \dqs_group[0].dq[6].dqi (
	.datain({dq_datain_6}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[6].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[6].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_8 \dqs_group[0].dq[7].dqi (
	.datain({dq_datain_7}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[0].dq[7].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[0].dq[7].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_9 \dqs_group[1].dq[0].dqi (
	.datain({dq_datain_8}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[0].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[0].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_10 \dqs_group[1].dq[1].dqi (
	.datain({dq_datain_9}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[1].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[1].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_11 \dqs_group[1].dq[2].dqi (
	.datain({dq_datain_10}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[2].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[2].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_12 \dqs_group[1].dq[3].dqi (
	.datain({dq_datain_11}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[3].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[3].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_13 \dqs_group[1].dq[4].dqi (
	.datain({dq_datain_12}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[4].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[4].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_14 \dqs_group[1].dq[5].dqi (
	.datain({dq_datain_13}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[5].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[5].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_15 \dqs_group[1].dq[6].dqi (
	.datain({dq_datain_14}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[6].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[6].dqi|auto_generated|input_cell_h[0]~q ));

altera_ddr_altddio_in_16 \dqs_group[1].dq[7].dqi (
	.datain({dq_datain_15}),
	.inclock(clk_3),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(\dqs_group[1].dq[7].dqi|auto_generated|input_latch_l[0]~q ),
	.input_cell_h_0(\dqs_group[1].dq[7].dqi|auto_generated|input_cell_h[0]~q ));

cycloneiii_ddio_out \dm[0].dm_ddio_out (
	.datainlo(wdp_dm_l_2x[0]),
	.datainhi(wdp_dm_h_2x[0]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dm_ddio_dataout_0),
	.dfflo(),
	.dffhi());
defparam \dm[0].dm_ddio_out .async_mode = "none";
defparam \dm[0].dm_ddio_out .power_up = "low";
defparam \dm[0].dm_ddio_out .sync_mode = "none";
defparam \dm[0].dm_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dm[1].dm_ddio_out (
	.datainlo(wdp_dm_l_2x[1]),
	.datainhi(wdp_dm_h_2x[1]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dm_ddio_dataout_1),
	.dfflo(),
	.dffhi());
defparam \dm[1].dm_ddio_out .async_mode = "none";
defparam \dm[1].dm_ddio_out .power_up = "low";
defparam \dm[1].dm_ddio_out .sync_mode = "none";
defparam \dm[1].dm_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[0].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[0]),
	.datainhi(wdp_wdata_h_2x[0]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_0),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[0].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[0].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[0].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[0].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[1].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[1]),
	.datainhi(wdp_wdata_h_2x[1]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_1),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[1].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[1].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[1].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[1].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[2].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[2]),
	.datainhi(wdp_wdata_h_2x[2]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_2),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[2].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[2].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[2].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[2].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[3].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[3]),
	.datainhi(wdp_wdata_h_2x[3]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_3),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[3].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[3].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[3].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[3].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[4].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[4]),
	.datainhi(wdp_wdata_h_2x[4]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_4),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[4].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[4].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[4].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[4].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[5].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[5]),
	.datainhi(wdp_wdata_h_2x[5]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_5),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[5].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[5].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[5].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[5].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[6].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[6]),
	.datainhi(wdp_wdata_h_2x[6]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_6),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[6].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[6].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[6].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[6].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[0].dq[7].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[7]),
	.datainhi(wdp_wdata_h_2x[7]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_7),
	.dfflo(),
	.dffhi());
defparam \dqs_group[0].dq[7].dq_ddio_out .async_mode = "none";
defparam \dqs_group[0].dq[7].dq_ddio_out .power_up = "low";
defparam \dqs_group[0].dq[7].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[0].dq[7].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[0].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[8]),
	.datainhi(wdp_wdata_h_2x[8]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_8),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[0].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[0].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[0].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[0].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[1].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[9]),
	.datainhi(wdp_wdata_h_2x[9]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_9),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[1].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[1].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[1].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[1].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[2].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[10]),
	.datainhi(wdp_wdata_h_2x[10]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_10),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[2].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[2].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[2].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[2].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[3].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[11]),
	.datainhi(wdp_wdata_h_2x[11]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_11),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[3].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[3].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[3].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[3].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[4].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[12]),
	.datainhi(wdp_wdata_h_2x[12]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_12),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[4].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[4].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[4].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[4].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[5].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[13]),
	.datainhi(wdp_wdata_h_2x[13]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_13),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[5].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[5].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[5].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[5].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[6].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[14]),
	.datainhi(wdp_wdata_h_2x[14]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_14),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[6].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[6].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[6].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[6].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs_group[1].dq[7].dq_ddio_out (
	.datainlo(wdp_wdata_l_2x[15]),
	.datainhi(wdp_wdata_h_2x[15]),
	.clkhi(write_clk_2x),
	.clklo(write_clk_2x),
	.muxsel(write_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dq_ddio_dataout_15),
	.dfflo(),
	.dffhi());
defparam \dqs_group[1].dq[7].dq_ddio_out .async_mode = "none";
defparam \dqs_group[1].dq[7].dq_ddio_out .power_up = "low";
defparam \dqs_group[1].dq[7].dq_ddio_out .sync_mode = "none";
defparam \dqs_group[1].dq[7].dq_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_out \dqs[0].dqs_ddio_out (
	.datainlo(gnd),
	.datainhi(wdp_wdqs_2x[0]),
	.clkhi(mem_clk_2x),
	.clklo(mem_clk_2x),
	.muxsel(mem_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dqs_ddio_dataout_0),
	.dfflo(),
	.dffhi());
defparam \dqs[0].dqs_ddio_out .async_mode = "none";
defparam \dqs[0].dqs_ddio_out .power_up = "low";
defparam \dqs[0].dqs_ddio_out .sync_mode = "none";
defparam \dqs[0].dqs_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_oe \dqs[0].dqsoe_ddio_oe (
	.oe(!wdp_wdqs_oe_2x[0]),
	.clk(mem_clk_2x),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(wdp_wdqs_oe_2x_r_0),
	.dfflo(),
	.dffhi());
defparam \dqs[0].dqsoe_ddio_oe .async_mode = "none";
defparam \dqs[0].dqsoe_ddio_oe .power_up = "low";
defparam \dqs[0].dqsoe_ddio_oe .sync_mode = "none";

cycloneiii_ddio_out \dqs[1].dqs_ddio_out (
	.datainlo(gnd),
	.datainhi(wdp_wdqs_2x[0]),
	.clkhi(mem_clk_2x),
	.clklo(mem_clk_2x),
	.muxsel(mem_clk_2x),
	.clk(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(dqs_ddio_dataout_1),
	.dfflo(),
	.dffhi());
defparam \dqs[1].dqs_ddio_out .async_mode = "none";
defparam \dqs[1].dqs_ddio_out .power_up = "low";
defparam \dqs[1].dqs_ddio_out .sync_mode = "none";
defparam \dqs[1].dqs_ddio_out .use_new_clocking_model = "true";

cycloneiii_ddio_oe \dqs[1].dqsoe_ddio_oe (
	.oe(!wdp_wdqs_oe_2x[0]),
	.clk(mem_clk_2x),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.dataout(wdp_wdqs_oe_2x_r_1),
	.dfflo(),
	.dffhi());
defparam \dqs[1].dqsoe_ddio_oe .async_mode = "none";
defparam \dqs[1].dqsoe_ddio_oe .power_up = "low";
defparam \dqs[1].dqsoe_ddio_oe .sync_mode = "none";

dffeas \wdp_wdata_oe_2x_r[0] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_0),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[0] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[0] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[1] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_1),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[1] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[1] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[2] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_2),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[2] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[2] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[3] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_3),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[3] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[3] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[4] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_4),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[4] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[4] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[5] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_5),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[5] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[5] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[6] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_6),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[6] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[6] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[7] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_7),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[7] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[7] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[8] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_8),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[8] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[8] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[9] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_9),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[9] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[9] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[10] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_10),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[10] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[10] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[11] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_11),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[11] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[11] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[12] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_12),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[12] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[12] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[13] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_13),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[13] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[13] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[14] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_14),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[14] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[14] .power_up = "low";

dffeas \wdp_wdata_oe_2x_r[15] (
	.clk(write_clk_2x),
	.d(wdp_wdata_oe_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_oe_2x_r_15),
	.prn(vcc));
defparam \wdp_wdata_oe_2x_r[15] .is_wysiwyg = "true";
defparam \wdp_wdata_oe_2x_r[15] .power_up = "low";

dffeas \dio_rdata_h_2x[0] (
	.clk(clk_3),
	.d(\rdata_p_ams[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_0),
	.prn(vcc));
defparam \dio_rdata_h_2x[0] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[0] .power_up = "low";

dffeas \dio_rdata_h_2x[1] (
	.clk(clk_3),
	.d(\rdata_p_ams[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_1),
	.prn(vcc));
defparam \dio_rdata_h_2x[1] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[1] .power_up = "low";

dffeas \dio_rdata_h_2x[2] (
	.clk(clk_3),
	.d(\rdata_p_ams[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_2),
	.prn(vcc));
defparam \dio_rdata_h_2x[2] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[2] .power_up = "low";

dffeas \dio_rdata_h_2x[3] (
	.clk(clk_3),
	.d(\rdata_p_ams[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_3),
	.prn(vcc));
defparam \dio_rdata_h_2x[3] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[3] .power_up = "low";

dffeas \dio_rdata_h_2x[4] (
	.clk(clk_3),
	.d(\rdata_p_ams[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_4),
	.prn(vcc));
defparam \dio_rdata_h_2x[4] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[4] .power_up = "low";

dffeas \dio_rdata_h_2x[5] (
	.clk(clk_3),
	.d(\rdata_p_ams[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_5),
	.prn(vcc));
defparam \dio_rdata_h_2x[5] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[5] .power_up = "low";

dffeas \dio_rdata_h_2x[6] (
	.clk(clk_3),
	.d(\rdata_p_ams[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_6),
	.prn(vcc));
defparam \dio_rdata_h_2x[6] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[6] .power_up = "low";

dffeas \dio_rdata_h_2x[7] (
	.clk(clk_3),
	.d(\rdata_p_ams[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_7),
	.prn(vcc));
defparam \dio_rdata_h_2x[7] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[7] .power_up = "low";

dffeas \dio_rdata_h_2x[8] (
	.clk(clk_3),
	.d(\rdata_p_ams[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_8),
	.prn(vcc));
defparam \dio_rdata_h_2x[8] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[8] .power_up = "low";

dffeas \dio_rdata_h_2x[9] (
	.clk(clk_3),
	.d(\rdata_p_ams[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_9),
	.prn(vcc));
defparam \dio_rdata_h_2x[9] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[9] .power_up = "low";

dffeas \dio_rdata_h_2x[10] (
	.clk(clk_3),
	.d(\rdata_p_ams[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_10),
	.prn(vcc));
defparam \dio_rdata_h_2x[10] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[10] .power_up = "low";

dffeas \dio_rdata_h_2x[11] (
	.clk(clk_3),
	.d(\rdata_p_ams[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_11),
	.prn(vcc));
defparam \dio_rdata_h_2x[11] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[11] .power_up = "low";

dffeas \dio_rdata_h_2x[12] (
	.clk(clk_3),
	.d(\rdata_p_ams[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_12),
	.prn(vcc));
defparam \dio_rdata_h_2x[12] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[12] .power_up = "low";

dffeas \dio_rdata_h_2x[13] (
	.clk(clk_3),
	.d(\rdata_p_ams[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_13),
	.prn(vcc));
defparam \dio_rdata_h_2x[13] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[13] .power_up = "low";

dffeas \dio_rdata_h_2x[14] (
	.clk(clk_3),
	.d(\rdata_p_ams[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_14),
	.prn(vcc));
defparam \dio_rdata_h_2x[14] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[14] .power_up = "low";

dffeas \dio_rdata_h_2x[15] (
	.clk(clk_3),
	.d(\rdata_p_ams[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_15),
	.prn(vcc));
defparam \dio_rdata_h_2x[15] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[15] .power_up = "low";

dffeas \dio_rdata_l_2x[0] (
	.clk(clk_3),
	.d(\rdata_n_ams[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_0),
	.prn(vcc));
defparam \dio_rdata_l_2x[0] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[0] .power_up = "low";

dffeas \dio_rdata_l_2x[1] (
	.clk(clk_3),
	.d(\rdata_n_ams[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_1),
	.prn(vcc));
defparam \dio_rdata_l_2x[1] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[1] .power_up = "low";

dffeas \dio_rdata_l_2x[2] (
	.clk(clk_3),
	.d(\rdata_n_ams[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_2),
	.prn(vcc));
defparam \dio_rdata_l_2x[2] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[2] .power_up = "low";

dffeas \dio_rdata_l_2x[3] (
	.clk(clk_3),
	.d(\rdata_n_ams[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_3),
	.prn(vcc));
defparam \dio_rdata_l_2x[3] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[3] .power_up = "low";

dffeas \dio_rdata_l_2x[4] (
	.clk(clk_3),
	.d(\rdata_n_ams[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_4),
	.prn(vcc));
defparam \dio_rdata_l_2x[4] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[4] .power_up = "low";

dffeas \dio_rdata_l_2x[5] (
	.clk(clk_3),
	.d(\rdata_n_ams[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_5),
	.prn(vcc));
defparam \dio_rdata_l_2x[5] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[5] .power_up = "low";

dffeas \dio_rdata_l_2x[6] (
	.clk(clk_3),
	.d(\rdata_n_ams[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_6),
	.prn(vcc));
defparam \dio_rdata_l_2x[6] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[6] .power_up = "low";

dffeas \dio_rdata_l_2x[7] (
	.clk(clk_3),
	.d(\rdata_n_ams[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_7),
	.prn(vcc));
defparam \dio_rdata_l_2x[7] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[7] .power_up = "low";

dffeas \dio_rdata_l_2x[8] (
	.clk(clk_3),
	.d(\rdata_n_ams[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_8),
	.prn(vcc));
defparam \dio_rdata_l_2x[8] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[8] .power_up = "low";

dffeas \dio_rdata_l_2x[9] (
	.clk(clk_3),
	.d(\rdata_n_ams[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_9),
	.prn(vcc));
defparam \dio_rdata_l_2x[9] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[9] .power_up = "low";

dffeas \dio_rdata_l_2x[10] (
	.clk(clk_3),
	.d(\rdata_n_ams[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_10),
	.prn(vcc));
defparam \dio_rdata_l_2x[10] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[10] .power_up = "low";

dffeas \dio_rdata_l_2x[11] (
	.clk(clk_3),
	.d(\rdata_n_ams[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_11),
	.prn(vcc));
defparam \dio_rdata_l_2x[11] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[11] .power_up = "low";

dffeas \dio_rdata_l_2x[12] (
	.clk(clk_3),
	.d(\rdata_n_ams[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_12),
	.prn(vcc));
defparam \dio_rdata_l_2x[12] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[12] .power_up = "low";

dffeas \dio_rdata_l_2x[13] (
	.clk(clk_3),
	.d(\rdata_n_ams[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_13),
	.prn(vcc));
defparam \dio_rdata_l_2x[13] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[13] .power_up = "low";

dffeas \dio_rdata_l_2x[14] (
	.clk(clk_3),
	.d(\rdata_n_ams[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_14),
	.prn(vcc));
defparam \dio_rdata_l_2x[14] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[14] .power_up = "low";

dffeas \dio_rdata_l_2x[15] (
	.clk(clk_3),
	.d(\rdata_n_ams[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_15),
	.prn(vcc));
defparam \dio_rdata_l_2x[15] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[15] .power_up = "low";

dffeas \rdata_p_ams[0] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[0].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[0]~q ),
	.prn(vcc));
defparam \rdata_p_ams[0] .is_wysiwyg = "true";
defparam \rdata_p_ams[0] .power_up = "low";

dffeas \rdata_p_ams[1] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[1].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[1]~q ),
	.prn(vcc));
defparam \rdata_p_ams[1] .is_wysiwyg = "true";
defparam \rdata_p_ams[1] .power_up = "low";

dffeas \rdata_p_ams[2] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[2].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[2]~q ),
	.prn(vcc));
defparam \rdata_p_ams[2] .is_wysiwyg = "true";
defparam \rdata_p_ams[2] .power_up = "low";

dffeas \rdata_p_ams[3] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[3].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[3]~q ),
	.prn(vcc));
defparam \rdata_p_ams[3] .is_wysiwyg = "true";
defparam \rdata_p_ams[3] .power_up = "low";

dffeas \rdata_p_ams[4] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[4].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[4]~q ),
	.prn(vcc));
defparam \rdata_p_ams[4] .is_wysiwyg = "true";
defparam \rdata_p_ams[4] .power_up = "low";

dffeas \rdata_p_ams[5] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[5].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[5]~q ),
	.prn(vcc));
defparam \rdata_p_ams[5] .is_wysiwyg = "true";
defparam \rdata_p_ams[5] .power_up = "low";

dffeas \rdata_p_ams[6] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[6].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[6]~q ),
	.prn(vcc));
defparam \rdata_p_ams[6] .is_wysiwyg = "true";
defparam \rdata_p_ams[6] .power_up = "low";

dffeas \rdata_p_ams[7] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[7].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[7]~q ),
	.prn(vcc));
defparam \rdata_p_ams[7] .is_wysiwyg = "true";
defparam \rdata_p_ams[7] .power_up = "low";

dffeas \rdata_p_ams[8] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[0].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[8]~q ),
	.prn(vcc));
defparam \rdata_p_ams[8] .is_wysiwyg = "true";
defparam \rdata_p_ams[8] .power_up = "low";

dffeas \rdata_p_ams[9] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[1].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[9]~q ),
	.prn(vcc));
defparam \rdata_p_ams[9] .is_wysiwyg = "true";
defparam \rdata_p_ams[9] .power_up = "low";

dffeas \rdata_p_ams[10] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[2].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[10]~q ),
	.prn(vcc));
defparam \rdata_p_ams[10] .is_wysiwyg = "true";
defparam \rdata_p_ams[10] .power_up = "low";

dffeas \rdata_p_ams[11] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[3].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[11]~q ),
	.prn(vcc));
defparam \rdata_p_ams[11] .is_wysiwyg = "true";
defparam \rdata_p_ams[11] .power_up = "low";

dffeas \rdata_p_ams[12] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[4].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[12]~q ),
	.prn(vcc));
defparam \rdata_p_ams[12] .is_wysiwyg = "true";
defparam \rdata_p_ams[12] .power_up = "low";

dffeas \rdata_p_ams[13] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[5].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[13]~q ),
	.prn(vcc));
defparam \rdata_p_ams[13] .is_wysiwyg = "true";
defparam \rdata_p_ams[13] .power_up = "low";

dffeas \rdata_p_ams[14] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[6].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[14]~q ),
	.prn(vcc));
defparam \rdata_p_ams[14] .is_wysiwyg = "true";
defparam \rdata_p_ams[14] .power_up = "low";

dffeas \rdata_p_ams[15] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[7].dqi|auto_generated|input_latch_l[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[15]~q ),
	.prn(vcc));
defparam \rdata_p_ams[15] .is_wysiwyg = "true";
defparam \rdata_p_ams[15] .power_up = "low";

dffeas \rdata_n_ams[0] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[0].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[0]~q ),
	.prn(vcc));
defparam \rdata_n_ams[0] .is_wysiwyg = "true";
defparam \rdata_n_ams[0] .power_up = "low";

dffeas \rdata_n_ams[1] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[1].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[1]~q ),
	.prn(vcc));
defparam \rdata_n_ams[1] .is_wysiwyg = "true";
defparam \rdata_n_ams[1] .power_up = "low";

dffeas \rdata_n_ams[2] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[2].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[2]~q ),
	.prn(vcc));
defparam \rdata_n_ams[2] .is_wysiwyg = "true";
defparam \rdata_n_ams[2] .power_up = "low";

dffeas \rdata_n_ams[3] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[3].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[3]~q ),
	.prn(vcc));
defparam \rdata_n_ams[3] .is_wysiwyg = "true";
defparam \rdata_n_ams[3] .power_up = "low";

dffeas \rdata_n_ams[4] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[4].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[4]~q ),
	.prn(vcc));
defparam \rdata_n_ams[4] .is_wysiwyg = "true";
defparam \rdata_n_ams[4] .power_up = "low";

dffeas \rdata_n_ams[5] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[5].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[5]~q ),
	.prn(vcc));
defparam \rdata_n_ams[5] .is_wysiwyg = "true";
defparam \rdata_n_ams[5] .power_up = "low";

dffeas \rdata_n_ams[6] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[6].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[6]~q ),
	.prn(vcc));
defparam \rdata_n_ams[6] .is_wysiwyg = "true";
defparam \rdata_n_ams[6] .power_up = "low";

dffeas \rdata_n_ams[7] (
	.clk(clk_3),
	.d(\dqs_group[0].dq[7].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[7]~q ),
	.prn(vcc));
defparam \rdata_n_ams[7] .is_wysiwyg = "true";
defparam \rdata_n_ams[7] .power_up = "low";

dffeas \rdata_n_ams[8] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[0].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[8]~q ),
	.prn(vcc));
defparam \rdata_n_ams[8] .is_wysiwyg = "true";
defparam \rdata_n_ams[8] .power_up = "low";

dffeas \rdata_n_ams[9] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[1].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[9]~q ),
	.prn(vcc));
defparam \rdata_n_ams[9] .is_wysiwyg = "true";
defparam \rdata_n_ams[9] .power_up = "low";

dffeas \rdata_n_ams[10] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[2].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[10]~q ),
	.prn(vcc));
defparam \rdata_n_ams[10] .is_wysiwyg = "true";
defparam \rdata_n_ams[10] .power_up = "low";

dffeas \rdata_n_ams[11] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[3].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[11]~q ),
	.prn(vcc));
defparam \rdata_n_ams[11] .is_wysiwyg = "true";
defparam \rdata_n_ams[11] .power_up = "low";

dffeas \rdata_n_ams[12] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[4].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[12]~q ),
	.prn(vcc));
defparam \rdata_n_ams[12] .is_wysiwyg = "true";
defparam \rdata_n_ams[12] .power_up = "low";

dffeas \rdata_n_ams[13] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[5].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[13]~q ),
	.prn(vcc));
defparam \rdata_n_ams[13] .is_wysiwyg = "true";
defparam \rdata_n_ams[13] .power_up = "low";

dffeas \rdata_n_ams[14] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[6].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[14]~q ),
	.prn(vcc));
defparam \rdata_n_ams[14] .is_wysiwyg = "true";
defparam \rdata_n_ams[14] .power_up = "low";

dffeas \rdata_n_ams[15] (
	.clk(clk_3),
	.d(\dqs_group[1].dq[7].dqi|auto_generated|input_cell_h[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[15]~q ),
	.prn(vcc));
defparam \rdata_n_ams[15] .is_wysiwyg = "true";
defparam \rdata_n_ams[15] .power_up = "low";

endmodule

module altera_ddr_altddio_in_1 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_2 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_1 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_1 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_3 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_2 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_2 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_4 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_3 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_3 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_5 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_4 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_4 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_6 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_5 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_5 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_7 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_6 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_6 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_8 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_7 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_7 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_9 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_8 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_8 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_10 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_9 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_9 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_11 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_10 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_10 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_12 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_11 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_11 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_13 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_12 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_12 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_14 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_13 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_13 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_15 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_14 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_14 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altddio_in_16 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_ddio_in_0fd_15 auto_generated(
	.datain({datain[0]}),
	.inclock(inclock),
	.ams_pipe_1(ams_pipe_1),
	.input_latch_l_0(input_latch_l_0),
	.input_cell_h_0(input_cell_h_0));

endmodule

module altera_ddr_ddio_in_0fd_15 (
	datain,
	inclock,
	ams_pipe_1,
	input_latch_l_0,
	input_cell_h_0)/* synthesis synthesis_greybox=1 */;
input 	[0:0] datain;
input 	inclock;
input 	ams_pipe_1;
output 	input_latch_l_0;
output 	input_cell_h_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \input_cell_l[0]~q ;


dffeas \input_latch_l[0] (
	.clk(inclock),
	.d(\input_cell_l[0]~q ),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_latch_l_0),
	.prn(vcc));
defparam \input_latch_l[0] .is_wysiwyg = "true";
defparam \input_latch_l[0] .power_up = "low";

dffeas \input_cell_h[0] (
	.clk(inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(input_cell_h_0),
	.prn(vcc));
defparam \input_cell_h[0] .is_wysiwyg = "true";
defparam \input_cell_h[0] .power_up = "low";

dffeas \input_cell_l[0] (
	.clk(!inclock),
	.d(datain[0]),
	.asdata(vcc),
	.clrn(ams_pipe_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\input_cell_l[0]~q ),
	.prn(vcc));
defparam \input_cell_l[0] .is_wysiwyg = "true";
defparam \input_cell_l[0] .power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_mimic (
	measure_clk,
	mimic_done_out1,
	reset_measure_clk_n,
	seq_mmc_start,
	mimic_value_captured1,
	mimic_data_in)/* synthesis synthesis_greybox=1 */;
input 	measure_clk;
output 	mimic_done_out1;
input 	reset_measure_clk_n;
input 	seq_mmc_start;
output 	mimic_value_captured1;
input 	mimic_data_in;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \shift_reg_counter[2]~q ;
wire \mimic_state.100~q ;
wire \start_edge_detected~0_combout ;
wire \Equal0~1_combout ;
wire \shift_reg_counter[2]~9_combout ;
wire \mimic_state.011~q ;
wire \mimic_state.010~q ;
wire \shift_reg_data_out[5]~q ;
wire \shift_reg_data_out[1]~q ;
wire \shift_reg_data_out~12_combout ;
wire \shift_reg_data_out~17_combout ;
wire \mimic_data_in_metastable[1]~q ;
wire \mimic_data_in_metastable[0]~q ;
wire \seq_mmc_start_metastable[0]~q ;
wire \seq_mmc_start_metastable[1]~q ;
wire \seq_mmc_start_metastable[2]~q ;
wire \Selector6~0_combout ;
wire \mimic_state.000~q ;
wire \shift_reg_counter[1]~8_combout ;
wire \Selector6~1_combout ;
wire \shift_reg_counter[0]~11_combout ;
wire \shift_reg_counter[0]~q ;
wire \shift_reg_counter[1]~10_combout ;
wire \shift_reg_counter[1]~q ;
wire \Equal0~2_combout ;
wire \shift_reg_counter[3]~12_combout ;
wire \shift_reg_counter[3]~q ;
wire \Equal0~0_combout ;
wire \Selector7~0_combout ;
wire \mimic_state.001~q ;
wire \Selector4~0_combout ;
wire \shift_reg_s_clr~0_combout ;
wire \shift_reg_s_clr~q ;
wire \shift_reg_data_out~14_combout ;
wire \Selector5~0_combout ;
wire \shift_reg_enable~q ;
wire \shift_reg_data_out[0]~13_combout ;
wire \shift_reg_data_out[4]~q ;
wire \shift_reg_data_out~15_combout ;
wire \shift_reg_data_out[3]~q ;
wire \shift_reg_data_out~16_combout ;
wire \shift_reg_data_out[2]~q ;
wire \mimic_value_captured~1_combout ;
wire \shift_reg_data_out~18_combout ;
wire \shift_reg_data_out[0]~q ;
wire \mimic_value_captured~2_combout ;
wire \shift_reg_counter[1]~13_combout ;
wire \mimic_value_captured~3_combout ;


dffeas \shift_reg_counter[2] (
	.clk(measure_clk),
	.d(\shift_reg_counter[2]~9_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[2]~q ),
	.prn(vcc));
defparam \shift_reg_counter[2] .is_wysiwyg = "true";
defparam \shift_reg_counter[2] .power_up = "low";

dffeas \mimic_state.100 (
	.clk(measure_clk),
	.d(\mimic_state.011~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.100~q ),
	.prn(vcc));
defparam \mimic_state.100 .is_wysiwyg = "true";
defparam \mimic_state.100 .power_up = "low";

cycloneiii_lcell_comb \start_edge_detected~0 (
	.dataa(\seq_mmc_start_metastable[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\seq_mmc_start_metastable[2]~q ),
	.cin(gnd),
	.combout(\start_edge_detected~0_combout ),
	.cout());
defparam \start_edge_detected~0 .lut_mask = 16'hAAFF;
defparam \start_edge_detected~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\shift_reg_counter[1]~q ),
	.datab(\shift_reg_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEEEE;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_counter[2]~9 (
	.dataa(\shift_reg_counter[2]~q ),
	.datab(\shift_reg_counter[1]~8_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\shift_reg_counter[2]~9_combout ),
	.cout());
defparam \shift_reg_counter[2]~9 .lut_mask = 16'h96FF;
defparam \shift_reg_counter[2]~9 .sum_lutc_input = "datac";

dffeas \mimic_state.011 (
	.clk(measure_clk),
	.d(\mimic_state.010~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.011~q ),
	.prn(vcc));
defparam \mimic_state.011 .is_wysiwyg = "true";
defparam \mimic_state.011 .power_up = "low";

dffeas \mimic_state.010 (
	.clk(measure_clk),
	.d(\shift_reg_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.010~q ),
	.prn(vcc));
defparam \mimic_state.010 .is_wysiwyg = "true";
defparam \mimic_state.010 .power_up = "low";

dffeas \shift_reg_data_out[5] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~12_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[5]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[5] .is_wysiwyg = "true";
defparam \shift_reg_data_out[5] .power_up = "low";

dffeas \shift_reg_data_out[1] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~17_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[1]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[1] .is_wysiwyg = "true";
defparam \shift_reg_data_out[1] .power_up = "low";

cycloneiii_lcell_comb \shift_reg_data_out~12 (
	.dataa(\shift_reg_data_out[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~12_combout ),
	.cout());
defparam \shift_reg_data_out~12 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_data_out~17 (
	.dataa(\shift_reg_data_out[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~17_combout ),
	.cout());
defparam \shift_reg_data_out~17 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~17 .sum_lutc_input = "datac";

dffeas \mimic_data_in_metastable[1] (
	.clk(measure_clk),
	.d(\mimic_data_in_metastable[0]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_data_in_metastable[1]~q ),
	.prn(vcc));
defparam \mimic_data_in_metastable[1] .is_wysiwyg = "true";
defparam \mimic_data_in_metastable[1] .power_up = "low";

dffeas \mimic_data_in_metastable[0] (
	.clk(measure_clk),
	.d(mimic_data_in),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_data_in_metastable[0]~q ),
	.prn(vcc));
defparam \mimic_data_in_metastable[0] .is_wysiwyg = "true";
defparam \mimic_data_in_metastable[0] .power_up = "low";

dffeas mimic_done_out(
	.clk(measure_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mimic_done_out1),
	.prn(vcc));
defparam mimic_done_out.is_wysiwyg = "true";
defparam mimic_done_out.power_up = "low";

dffeas mimic_value_captured(
	.clk(measure_clk),
	.d(\mimic_value_captured~3_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mimic_value_captured1),
	.prn(vcc));
defparam mimic_value_captured.is_wysiwyg = "true";
defparam mimic_value_captured.power_up = "low";

dffeas \seq_mmc_start_metastable[0] (
	.clk(measure_clk),
	.d(seq_mmc_start),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[0]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[0] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[0] .power_up = "low";

dffeas \seq_mmc_start_metastable[1] (
	.clk(measure_clk),
	.d(\seq_mmc_start_metastable[0]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[1]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[1] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[1] .power_up = "low";

dffeas \seq_mmc_start_metastable[2] (
	.clk(measure_clk),
	.d(\seq_mmc_start_metastable[1]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[2]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[2] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[2] .power_up = "low";

cycloneiii_lcell_comb \Selector6~0 (
	.dataa(\mimic_state.100~q ),
	.datab(\seq_mmc_start_metastable[2]~q ),
	.datac(\seq_mmc_start_metastable[1]~q ),
	.datad(\mimic_state.000~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hFFF7;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \mimic_state.000 (
	.clk(measure_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.000~q ),
	.prn(vcc));
defparam \mimic_state.000 .is_wysiwyg = "true";
defparam \mimic_state.000 .power_up = "low";

cycloneiii_lcell_comb \shift_reg_counter[1]~8 (
	.dataa(\Equal0~0_combout ),
	.datab(\mimic_state.000~q ),
	.datac(gnd),
	.datad(\mimic_state.001~q ),
	.cin(gnd),
	.combout(\shift_reg_counter[1]~8_combout ),
	.cout());
defparam \shift_reg_counter[1]~8 .lut_mask = 16'hAACC;
defparam \shift_reg_counter[1]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~1 (
	.dataa(\seq_mmc_start_metastable[2]~q ),
	.datab(gnd),
	.datac(\seq_mmc_start_metastable[1]~q ),
	.datad(\mimic_state.000~q ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hAFFF;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_counter[0]~11 (
	.dataa(\shift_reg_counter[0]~q ),
	.datab(\shift_reg_counter[1]~8_combout ),
	.datac(gnd),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\shift_reg_counter[0]~11_combout ),
	.cout());
defparam \shift_reg_counter[0]~11 .lut_mask = 16'h66FF;
defparam \shift_reg_counter[0]~11 .sum_lutc_input = "datac";

dffeas \shift_reg_counter[0] (
	.clk(measure_clk),
	.d(\shift_reg_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[0]~q ),
	.prn(vcc));
defparam \shift_reg_counter[0] .is_wysiwyg = "true";
defparam \shift_reg_counter[0] .power_up = "low";

cycloneiii_lcell_comb \shift_reg_counter[1]~10 (
	.dataa(\shift_reg_counter[1]~q ),
	.datab(\shift_reg_counter[1]~8_combout ),
	.datac(\shift_reg_counter[0]~q ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\shift_reg_counter[1]~10_combout ),
	.cout());
defparam \shift_reg_counter[1]~10 .lut_mask = 16'h96FF;
defparam \shift_reg_counter[1]~10 .sum_lutc_input = "datac";

dffeas \shift_reg_counter[1] (
	.clk(measure_clk),
	.d(\shift_reg_counter[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[1]~q ),
	.prn(vcc));
defparam \shift_reg_counter[1] .is_wysiwyg = "true";
defparam \shift_reg_counter[1] .power_up = "low";

cycloneiii_lcell_comb \Equal0~2 (
	.dataa(\shift_reg_counter[2]~q ),
	.datab(\shift_reg_counter[1]~q ),
	.datac(\shift_reg_counter[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFEFE;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_counter[3]~12 (
	.dataa(\shift_reg_counter[3]~q ),
	.datab(\shift_reg_counter[1]~8_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\shift_reg_counter[3]~12_combout ),
	.cout());
defparam \shift_reg_counter[3]~12 .lut_mask = 16'h96FF;
defparam \shift_reg_counter[3]~12 .sum_lutc_input = "datac";

dffeas \shift_reg_counter[3] (
	.clk(measure_clk),
	.d(\shift_reg_counter[3]~12_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[3]~q ),
	.prn(vcc));
defparam \shift_reg_counter[3] .is_wysiwyg = "true";
defparam \shift_reg_counter[3] .power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\shift_reg_counter[2]~q ),
	.datab(\shift_reg_counter[1]~q ),
	.datac(\shift_reg_counter[0]~q ),
	.datad(\shift_reg_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(\start_edge_detected~0_combout ),
	.datab(\mimic_state.001~q ),
	.datac(\mimic_state.000~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEFFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \mimic_state.001 (
	.clk(measure_clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.001~q ),
	.prn(vcc));
defparam \mimic_state.001 .is_wysiwyg = "true";
defparam \mimic_state.001 .power_up = "low";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\mimic_state.000~q ),
	.datab(\mimic_state.001~q ),
	.datac(mimic_done_out1),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFFB8;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_s_clr~0 (
	.dataa(\shift_reg_s_clr~q ),
	.datab(\seq_mmc_start_metastable[2]~q ),
	.datac(\seq_mmc_start_metastable[1]~q ),
	.datad(\mimic_state.000~q ),
	.cin(gnd),
	.combout(\shift_reg_s_clr~0_combout ),
	.cout());
defparam \shift_reg_s_clr~0 .lut_mask = 16'hAFCF;
defparam \shift_reg_s_clr~0 .sum_lutc_input = "datac";

dffeas shift_reg_s_clr(
	.clk(measure_clk),
	.d(\shift_reg_s_clr~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_s_clr~q ),
	.prn(vcc));
defparam shift_reg_s_clr.is_wysiwyg = "true";
defparam shift_reg_s_clr.power_up = "low";

cycloneiii_lcell_comb \shift_reg_data_out~14 (
	.dataa(\shift_reg_data_out[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~14_combout ),
	.cout());
defparam \shift_reg_data_out~14 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\shift_reg_enable~q ),
	.datab(\mimic_state.000~q ),
	.datac(\Equal0~0_combout ),
	.datad(\mimic_state.001~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hBFFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas shift_reg_enable(
	.clk(measure_clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_enable~q ),
	.prn(vcc));
defparam shift_reg_enable.is_wysiwyg = "true";
defparam shift_reg_enable.power_up = "low";

cycloneiii_lcell_comb \shift_reg_data_out[0]~13 (
	.dataa(\shift_reg_s_clr~q ),
	.datab(\shift_reg_enable~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\shift_reg_data_out[0]~13_combout ),
	.cout());
defparam \shift_reg_data_out[0]~13 .lut_mask = 16'hEEEE;
defparam \shift_reg_data_out[0]~13 .sum_lutc_input = "datac";

dffeas \shift_reg_data_out[4] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~14_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[4]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[4] .is_wysiwyg = "true";
defparam \shift_reg_data_out[4] .power_up = "low";

cycloneiii_lcell_comb \shift_reg_data_out~15 (
	.dataa(\shift_reg_data_out[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~15_combout ),
	.cout());
defparam \shift_reg_data_out~15 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~15 .sum_lutc_input = "datac";

dffeas \shift_reg_data_out[3] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~15_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[3]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[3] .is_wysiwyg = "true";
defparam \shift_reg_data_out[3] .power_up = "low";

cycloneiii_lcell_comb \shift_reg_data_out~16 (
	.dataa(\shift_reg_data_out[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~16_combout ),
	.cout());
defparam \shift_reg_data_out~16 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~16 .sum_lutc_input = "datac";

dffeas \shift_reg_data_out[2] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~16_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[2]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[2] .is_wysiwyg = "true";
defparam \shift_reg_data_out[2] .power_up = "low";

cycloneiii_lcell_comb \mimic_value_captured~1 (
	.dataa(\shift_reg_data_out[5]~q ),
	.datab(\shift_reg_data_out[4]~q ),
	.datac(\shift_reg_data_out[3]~q ),
	.datad(\shift_reg_data_out[2]~q ),
	.cin(gnd),
	.combout(\mimic_value_captured~1_combout ),
	.cout());
defparam \mimic_value_captured~1 .lut_mask = 16'hFFFE;
defparam \mimic_value_captured~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_data_out~18 (
	.dataa(\mimic_data_in_metastable[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\shift_reg_s_clr~q ),
	.cin(gnd),
	.combout(\shift_reg_data_out~18_combout ),
	.cout());
defparam \shift_reg_data_out~18 .lut_mask = 16'hAAFF;
defparam \shift_reg_data_out~18 .sum_lutc_input = "datac";

dffeas \shift_reg_data_out[0] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~18_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~13_combout ),
	.q(\shift_reg_data_out[0]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[0] .is_wysiwyg = "true";
defparam \shift_reg_data_out[0] .power_up = "low";

cycloneiii_lcell_comb \mimic_value_captured~2 (
	.dataa(\shift_reg_data_out[1]~q ),
	.datab(\shift_reg_data_out[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mimic_value_captured~2_combout ),
	.cout());
defparam \mimic_value_captured~2 .lut_mask = 16'hEEEE;
defparam \mimic_value_captured~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \shift_reg_counter[1]~13 (
	.dataa(\mimic_state.001~q ),
	.datab(\Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\shift_reg_counter[1]~13_combout ),
	.cout());
defparam \shift_reg_counter[1]~13 .lut_mask = 16'hEEEE;
defparam \shift_reg_counter[1]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mimic_value_captured~3 (
	.dataa(\mimic_value_captured~1_combout ),
	.datab(\mimic_value_captured~2_combout ),
	.datac(mimic_value_captured1),
	.datad(\shift_reg_counter[1]~13_combout ),
	.cin(gnd),
	.combout(\mimic_value_captured~3_combout ),
	.cout());
defparam \mimic_value_captured~3 .lut_mask = 16'hFAFC;
defparam \mimic_value_captured~3 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_rdata_valid (
	clk_1,
	ctl_rdata_valid_0,
	ctl_init_success,
	reset_phy_clk_1x_n,
	rd_addr_0,
	rd_ram_rd_addr_1,
	rd_ram_rd_addr_2,
	rd_ram_rd_addr_3,
	seq_rdv_doing_rd_0,
	seq_rdv_doing_rd_1,
	control_doing_rd_0,
	seq_rdata_valid_lat_dec,
	Add2,
	seq_rdata_valid_0)/* synthesis synthesis_greybox=1 */;
input 	clk_1;
output 	ctl_rdata_valid_0;
input 	ctl_init_success;
input 	reset_phy_clk_1x_n;
output 	rd_addr_0;
input 	rd_ram_rd_addr_1;
input 	rd_ram_rd_addr_2;
input 	rd_ram_rd_addr_3;
input 	seq_rdv_doing_rd_0;
input 	seq_rdv_doing_rd_1;
input 	control_doing_rd_0;
input 	seq_rdata_valid_lat_dec;
input 	Add2;
output 	seq_rdata_valid_0;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \altsyncram_component|auto_generated|q_b[0] ;
wire \wr_addr[1]~q ;
wire \wr_addr[2]~q ;
wire \wr_addr[3]~q ;
wire \wr_addr[4]~q ;
wire \wr_addr[1]~11 ;
wire \wr_addr[1]~10_combout ;
wire \wr_addr[2]~13 ;
wire \wr_addr[2]~12_combout ;
wire \wr_addr[3]~15 ;
wire \wr_addr[3]~14_combout ;
wire \wr_addr[4]~16_combout ;
wire \WideOr0~combout ;
wire \wr_addr[0]~q ;
wire \rd_addr[4]~q ;
wire \seq_rdata_valid_lat_dec_1t~q ;
wire \wr_addr[0]~9_combout ;
wire \always3~0_combout ;
wire \rd_addr[4]~5_combout ;
wire \wr_addr[0]~_wirecell_combout ;
wire \wr_addr[1]~_wirecell_combout ;
wire \wr_addr[2]~_wirecell_combout ;
wire \wr_addr[4]~_wirecell_combout ;
wire \ctl_rdata_valid~0_combout ;
wire \rd_addr[0]~6_combout ;


altera_ddr_altsyncram_1 altsyncram_component(
	.clock0(clk_1),
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,\altsyncram_component|auto_generated|q_b[0] }),
	.address_a({\wr_addr[4]~_wirecell_combout ,\wr_addr[3]~q ,\wr_addr[2]~_wirecell_combout ,\wr_addr[1]~_wirecell_combout ,\wr_addr[0]~_wirecell_combout }),
	.address_b({\rd_addr[4]~q ,rd_ram_rd_addr_3,rd_ram_rd_addr_2,rd_ram_rd_addr_1,rd_addr_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\WideOr0~combout }));

dffeas \wr_addr[1] (
	.clk(clk_1),
	.d(\wr_addr[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\wr_addr[1]~q ),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

dffeas \wr_addr[2] (
	.clk(clk_1),
	.d(\wr_addr[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\wr_addr[2]~q ),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

dffeas \wr_addr[3] (
	.clk(clk_1),
	.d(\wr_addr[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\wr_addr[3]~q ),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

dffeas \wr_addr[4] (
	.clk(clk_1),
	.d(\wr_addr[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\wr_addr[4]~q ),
	.prn(vcc));
defparam \wr_addr[4] .is_wysiwyg = "true";
defparam \wr_addr[4] .power_up = "low";

cycloneiii_lcell_comb \wr_addr[1]~10 (
	.dataa(\wr_addr[0]~q ),
	.datab(\wr_addr[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\wr_addr[1]~10_combout ),
	.cout(\wr_addr[1]~11 ));
defparam \wr_addr[1]~10 .lut_mask = 16'h6677;
defparam \wr_addr[1]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wr_addr[2]~12 (
	.dataa(\wr_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\wr_addr[1]~11 ),
	.combout(\wr_addr[2]~12_combout ),
	.cout(\wr_addr[2]~13 ));
defparam \wr_addr[2]~12 .lut_mask = 16'h5AAF;
defparam \wr_addr[2]~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \wr_addr[3]~14 (
	.dataa(\wr_addr[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\wr_addr[2]~13 ),
	.combout(\wr_addr[3]~14_combout ),
	.cout(\wr_addr[3]~15 ));
defparam \wr_addr[3]~14 .lut_mask = 16'h5AAF;
defparam \wr_addr[3]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \wr_addr[4]~16 (
	.dataa(\wr_addr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\wr_addr[3]~15 ),
	.combout(\wr_addr[4]~16_combout ),
	.cout());
defparam \wr_addr[4]~16 .lut_mask = 16'h5A5A;
defparam \wr_addr[4]~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb WideOr0(
	.dataa(seq_rdv_doing_rd_0),
	.datab(seq_rdv_doing_rd_1),
	.datac(ctl_init_success),
	.datad(control_doing_rd_0),
	.cin(gnd),
	.combout(\WideOr0~combout ),
	.cout());
defparam WideOr0.lut_mask = 16'hFFFE;
defparam WideOr0.sum_lutc_input = "datac";

dffeas \wr_addr[0] (
	.clk(clk_1),
	.d(\wr_addr[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_addr[0]~q ),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

dffeas \rd_addr[4] (
	.clk(clk_1),
	.d(\rd_addr[4]~5_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr[4]~q ),
	.prn(vcc));
defparam \rd_addr[4] .is_wysiwyg = "true";
defparam \rd_addr[4] .power_up = "low";

dffeas seq_rdata_valid_lat_dec_1t(
	.clk(clk_1),
	.d(seq_rdata_valid_lat_dec),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_rdata_valid_lat_dec_1t~q ),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec_1t.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec_1t.power_up = "low";

cycloneiii_lcell_comb \wr_addr[0]~9 (
	.dataa(seq_rdata_valid_lat_dec),
	.datab(gnd),
	.datac(\seq_rdata_valid_lat_dec_1t~q ),
	.datad(\wr_addr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr[0]~9_combout ),
	.cout());
defparam \wr_addr[0]~9 .lut_mask = 16'hA55A;
defparam \wr_addr[0]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \always3~0 (
	.dataa(seq_rdata_valid_lat_dec),
	.datab(gnd),
	.datac(gnd),
	.datad(\seq_rdata_valid_lat_dec_1t~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'hFF55;
defparam \always3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_addr[4]~5 (
	.dataa(\rd_addr[4]~q ),
	.datab(rd_ram_rd_addr_2),
	.datac(rd_ram_rd_addr_3),
	.datad(Add2),
	.cin(gnd),
	.combout(\rd_addr[4]~5_combout ),
	.cout());
defparam \rd_addr[4]~5 .lut_mask = 16'h6996;
defparam \rd_addr[4]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wr_addr[0]~_wirecell (
	.dataa(\wr_addr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_addr[0]~_wirecell_combout ),
	.cout());
defparam \wr_addr[0]~_wirecell .lut_mask = 16'h5555;
defparam \wr_addr[0]~_wirecell .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wr_addr[1]~_wirecell (
	.dataa(\wr_addr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_addr[1]~_wirecell_combout ),
	.cout());
defparam \wr_addr[1]~_wirecell .lut_mask = 16'h5555;
defparam \wr_addr[1]~_wirecell .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wr_addr[2]~_wirecell (
	.dataa(\wr_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_addr[2]~_wirecell_combout ),
	.cout());
defparam \wr_addr[2]~_wirecell .lut_mask = 16'h5555;
defparam \wr_addr[2]~_wirecell .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wr_addr[4]~_wirecell (
	.dataa(\wr_addr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_addr[4]~_wirecell_combout ),
	.cout());
defparam \wr_addr[4]~_wirecell .lut_mask = 16'h5555;
defparam \wr_addr[4]~_wirecell .sum_lutc_input = "datac";

dffeas \ctl_rdata_valid[0] (
	.clk(clk_1),
	.d(\ctl_rdata_valid~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_rdata_valid_0),
	.prn(vcc));
defparam \ctl_rdata_valid[0] .is_wysiwyg = "true";
defparam \ctl_rdata_valid[0] .power_up = "low";

dffeas \rd_addr[0] (
	.clk(clk_1),
	.d(\rd_addr[0]~6_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_addr_0),
	.prn(vcc));
defparam \rd_addr[0] .is_wysiwyg = "true";
defparam \rd_addr[0] .power_up = "low";

dffeas \seq_rdata_valid[0] (
	.clk(clk_1),
	.d(\altsyncram_component|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_0),
	.prn(vcc));
defparam \seq_rdata_valid[0] .is_wysiwyg = "true";
defparam \seq_rdata_valid[0] .power_up = "low";

cycloneiii_lcell_comb \ctl_rdata_valid~0 (
	.dataa(ctl_init_success),
	.datab(\altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ctl_rdata_valid~0_combout ),
	.cout());
defparam \ctl_rdata_valid~0 .lut_mask = 16'hEEEE;
defparam \ctl_rdata_valid~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_addr[0]~6 (
	.dataa(rd_addr_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_addr[0]~6_combout ),
	.cout());
defparam \rd_addr[0]~6 .lut_mask = 16'h5555;
defparam \rd_addr[0]~6 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altsyncram_1 (
	clock0,
	q_b,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[31:0] q_b;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	[31:0] data_a;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altsyncram_2ni1 auto_generated(
	.clock0(clock0),
	.q_b({q_b[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[0]}));

endmodule

module altera_ddr_altsyncram_2ni1 (
	clock0,
	q_b,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=1 */;
input 	clock0;
output 	[0:0] q_b;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	[0:0] data_a;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_rdata_valid:rdv_pipe|altsyncram:altsyncram_component|altsyncram_2ni1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 1;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 1;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_read_dp (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk_1,
	clk_3,
	reset_phy_clk_1x_n,
	rd_addr_0,
	rd_ram_rd_addr_1,
	rd_ram_rd_addr_2,
	rd_ram_rd_addr_3,
	reset_resync_clk_2x_n,
	dio_rdata_h_2x,
	dio_rdata_l_2x,
	Add2)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_24;
output 	q_b_25;
output 	q_b_26;
output 	q_b_27;
output 	q_b_28;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
input 	clk_1;
input 	clk_3;
input 	reset_phy_clk_1x_n;
input 	rd_addr_0;
output 	rd_ram_rd_addr_1;
output 	rd_ram_rd_addr_2;
output 	rd_ram_rd_addr_3;
input 	reset_resync_clk_2x_n;
input 	[15:0] dio_rdata_h_2x;
input 	[15:0] dio_rdata_l_2x;
output 	Add2;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \resync_pipeline_gen.pipeline_delay[1][0]~q ;
wire \rd_ram_wr_addr[0]~q ;
wire \rd_ram_wr_addr[1]~q ;
wire \rd_ram_wr_addr[2]~q ;
wire \rd_ram_wr_addr[3]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][1]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][2]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][3]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][4]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][5]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][6]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][7]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][16]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][17]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][18]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][19]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][20]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][21]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][22]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][23]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][8]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][9]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][10]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][11]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][12]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][13]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][14]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][15]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][24]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][25]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][26]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][27]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][28]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][29]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][30]~q ;
wire \resync_pipeline_gen.pipeline_delay[1][31]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][0]~q ;
wire \rd_ram_wr_addr[1]~8_combout ;
wire \rd_ram_wr_addr[2]~9_combout ;
wire \rd_ram_wr_addr[3]~10_combout ;
wire \resync_pipeline_gen.pipeline_delay[0][1]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][2]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][3]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][4]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][5]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][6]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][7]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][16]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][17]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][18]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][19]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][20]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][21]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][22]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][23]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][8]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][9]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][10]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][11]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][12]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][13]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][14]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][15]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][24]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][25]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][26]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][27]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][28]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][29]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][30]~q ;
wire \resync_pipeline_gen.pipeline_delay[0][31]~q ;
wire \rd_ram_wr_addr[0]~11_combout ;
wire \rd_ram_wr_addr[1]~_wirecell_combout ;
wire \rd_ram_wr_addr[2]~_wirecell_combout ;
wire \rd_ram_rd_addr[1]~8_combout ;
wire \rd_ram_rd_addr[2]~9_combout ;
wire \rd_ram_rd_addr[3]~10_combout ;


altera_ddr_altsyncram_2 \full_rate_ram_gen.altsyncram_component (
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clock1(clk_1),
	.clock0(clk_3),
	.data_a({\resync_pipeline_gen.pipeline_delay[1][31]~q ,\resync_pipeline_gen.pipeline_delay[1][30]~q ,\resync_pipeline_gen.pipeline_delay[1][29]~q ,\resync_pipeline_gen.pipeline_delay[1][28]~q ,\resync_pipeline_gen.pipeline_delay[1][27]~q ,
\resync_pipeline_gen.pipeline_delay[1][26]~q ,\resync_pipeline_gen.pipeline_delay[1][25]~q ,\resync_pipeline_gen.pipeline_delay[1][24]~q ,\resync_pipeline_gen.pipeline_delay[1][23]~q ,\resync_pipeline_gen.pipeline_delay[1][22]~q ,
\resync_pipeline_gen.pipeline_delay[1][21]~q ,\resync_pipeline_gen.pipeline_delay[1][20]~q ,\resync_pipeline_gen.pipeline_delay[1][19]~q ,\resync_pipeline_gen.pipeline_delay[1][18]~q ,\resync_pipeline_gen.pipeline_delay[1][17]~q ,
\resync_pipeline_gen.pipeline_delay[1][16]~q ,\resync_pipeline_gen.pipeline_delay[1][15]~q ,\resync_pipeline_gen.pipeline_delay[1][14]~q ,\resync_pipeline_gen.pipeline_delay[1][13]~q ,\resync_pipeline_gen.pipeline_delay[1][12]~q ,
\resync_pipeline_gen.pipeline_delay[1][11]~q ,\resync_pipeline_gen.pipeline_delay[1][10]~q ,\resync_pipeline_gen.pipeline_delay[1][9]~q ,\resync_pipeline_gen.pipeline_delay[1][8]~q ,\resync_pipeline_gen.pipeline_delay[1][7]~q ,
\resync_pipeline_gen.pipeline_delay[1][6]~q ,\resync_pipeline_gen.pipeline_delay[1][5]~q ,\resync_pipeline_gen.pipeline_delay[1][4]~q ,\resync_pipeline_gen.pipeline_delay[1][3]~q ,\resync_pipeline_gen.pipeline_delay[1][2]~q ,
\resync_pipeline_gen.pipeline_delay[1][1]~q ,\resync_pipeline_gen.pipeline_delay[1][0]~q }),
	.address_a({gnd,\rd_ram_wr_addr[3]~q ,\rd_ram_wr_addr[2]~_wirecell_combout ,\rd_ram_wr_addr[1]~_wirecell_combout ,\rd_ram_wr_addr[0]~q }),
	.address_b({gnd,rd_ram_rd_addr_3,rd_ram_rd_addr_2,rd_ram_rd_addr_1,rd_addr_0}));

dffeas \resync_pipeline_gen.pipeline_delay[1][0] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][0]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][0] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][0] .power_up = "low";

dffeas \rd_ram_wr_addr[0] (
	.clk(clk_3),
	.d(\rd_ram_wr_addr[0]~11_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[0]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[0] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[0] .power_up = "low";

dffeas \rd_ram_wr_addr[1] (
	.clk(clk_3),
	.d(\rd_ram_wr_addr[1]~8_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[1]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[1] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[1] .power_up = "low";

dffeas \rd_ram_wr_addr[2] (
	.clk(clk_3),
	.d(\rd_ram_wr_addr[2]~9_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[2]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[2] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[2] .power_up = "low";

dffeas \rd_ram_wr_addr[3] (
	.clk(clk_3),
	.d(\rd_ram_wr_addr[3]~10_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[3]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[3] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[3] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][1] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][1]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][1] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][1] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][2] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][2]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][2] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][2] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][3] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][3]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][3] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][3] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][4] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][4]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][4] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][4] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][5] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][5]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][5] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][5] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][6] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][6]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][6] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][6] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][7] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][7]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][7] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][7] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][16] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][16]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][16] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][16] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][17] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][17]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][17] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][17] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][18] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][18]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][18] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][18] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][19] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][19]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][19] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][19] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][20] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][20]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][20] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][20] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][21] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][21]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][21] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][21] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][22] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][22]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][22] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][22] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][23] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][23]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][23] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][23] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][8] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][8]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][8] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][8] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][9] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][9]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][9] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][9] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][10] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][10]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][10] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][10] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][11] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][11]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][11] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][11] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][12] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][12]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][12] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][12] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][13] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][13]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][13] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][13] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][14] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][14]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][14] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][14] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][15] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][15]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][15] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][15] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][24] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][24]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][24] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][24] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][25] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][25]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][25] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][25] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][26] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][26]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][26] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][26] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][27] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][27]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][27] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][27] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][28] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][28]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][28] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][28] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][29] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][29]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][29] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][29] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][30] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][30]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][30] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][30] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[1][31] (
	.clk(clk_3),
	.d(\resync_pipeline_gen.pipeline_delay[0][31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[1][31]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[1][31] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[1][31] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][0] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][0]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][0] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][0] .power_up = "low";

cycloneiii_lcell_comb \rd_ram_wr_addr[1]~8 (
	.dataa(\rd_ram_wr_addr[0]~q ),
	.datab(\rd_ram_wr_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[1]~8_combout ),
	.cout());
defparam \rd_ram_wr_addr[1]~8 .lut_mask = 16'h6666;
defparam \rd_ram_wr_addr[1]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_wr_addr[2]~9 (
	.dataa(\rd_ram_wr_addr[0]~q ),
	.datab(gnd),
	.datac(\rd_ram_wr_addr[1]~q ),
	.datad(\rd_ram_wr_addr[2]~q ),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[2]~9_combout ),
	.cout());
defparam \rd_ram_wr_addr[2]~9 .lut_mask = 16'hA55A;
defparam \rd_ram_wr_addr[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_wr_addr[3]~10 (
	.dataa(\rd_ram_wr_addr[3]~q ),
	.datab(\rd_ram_wr_addr[1]~q ),
	.datac(\rd_ram_wr_addr[2]~q ),
	.datad(\rd_ram_wr_addr[0]~q ),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[3]~10_combout ),
	.cout());
defparam \rd_ram_wr_addr[3]~10 .lut_mask = 16'h6996;
defparam \rd_ram_wr_addr[3]~10 .sum_lutc_input = "datac";

dffeas \resync_pipeline_gen.pipeline_delay[0][1] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][1]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][1] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][1] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][2] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][2]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][2] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][2] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][3] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][3]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][3] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][3] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][4] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][4]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][4] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][4] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][5] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][5]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][5] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][5] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][6] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][6]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][6] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][6] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][7] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][7]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][7] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][7] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][16] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][16]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][16] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][16] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][17] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][17]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][17] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][17] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][18] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][18]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][18] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][18] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][19] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][19]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][19] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][19] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][20] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][20]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][20] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][20] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][21] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][21]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][21] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][21] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][22] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][22]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][22] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][22] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][23] (
	.clk(clk_3),
	.d(dio_rdata_h_2x[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][23]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][23] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][23] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][8] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][8]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][8] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][8] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][9] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][9]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][9] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][9] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][10] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][10]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][10] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][10] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][11] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][11]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][11] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][11] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][12] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][12]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][12] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][12] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][13] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][13]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][13] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][13] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][14] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][14]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][14] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][14] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][15] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][15]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][15] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][15] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][24] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][24]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][24] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][24] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][25] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][25]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][25] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][25] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][26] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][26]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][26] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][26] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][27] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][27]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][27] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][27] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][28] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][28]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][28] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][28] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][29] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][29]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][29] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][29] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][30] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][30]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][30] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][30] .power_up = "low";

dffeas \resync_pipeline_gen.pipeline_delay[0][31] (
	.clk(clk_3),
	.d(dio_rdata_l_2x[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\resync_pipeline_gen.pipeline_delay[0][31]~q ),
	.prn(vcc));
defparam \resync_pipeline_gen.pipeline_delay[0][31] .is_wysiwyg = "true";
defparam \resync_pipeline_gen.pipeline_delay[0][31] .power_up = "low";

cycloneiii_lcell_comb \rd_ram_wr_addr[0]~11 (
	.dataa(\rd_ram_wr_addr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[0]~11_combout ),
	.cout());
defparam \rd_ram_wr_addr[0]~11 .lut_mask = 16'h5555;
defparam \rd_ram_wr_addr[0]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_wr_addr[1]~_wirecell (
	.dataa(\rd_ram_wr_addr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[1]~_wirecell_combout ),
	.cout());
defparam \rd_ram_wr_addr[1]~_wirecell .lut_mask = 16'h5555;
defparam \rd_ram_wr_addr[1]~_wirecell .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_wr_addr[2]~_wirecell (
	.dataa(\rd_ram_wr_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_ram_wr_addr[2]~_wirecell_combout ),
	.cout());
defparam \rd_ram_wr_addr[2]~_wirecell .lut_mask = 16'h5555;
defparam \rd_ram_wr_addr[2]~_wirecell .sum_lutc_input = "datac";

dffeas \rd_ram_rd_addr[1] (
	.clk(clk_1),
	.d(\rd_ram_rd_addr[1]~8_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_ram_rd_addr_1),
	.prn(vcc));
defparam \rd_ram_rd_addr[1] .is_wysiwyg = "true";
defparam \rd_ram_rd_addr[1] .power_up = "low";

dffeas \rd_ram_rd_addr[2] (
	.clk(clk_1),
	.d(\rd_ram_rd_addr[2]~9_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_ram_rd_addr_2),
	.prn(vcc));
defparam \rd_ram_rd_addr[2] .is_wysiwyg = "true";
defparam \rd_ram_rd_addr[2] .power_up = "low";

dffeas \rd_ram_rd_addr[3] (
	.clk(clk_1),
	.d(\rd_ram_rd_addr[3]~10_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_ram_rd_addr_3),
	.prn(vcc));
defparam \rd_ram_rd_addr[3] .is_wysiwyg = "true";
defparam \rd_ram_rd_addr[3] .power_up = "low";

cycloneiii_lcell_comb \Add2~0 (
	.dataa(rd_addr_0),
	.datab(rd_ram_rd_addr_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Add2),
	.cout());
defparam \Add2~0 .lut_mask = 16'hEEEE;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_rd_addr[1]~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(rd_addr_0),
	.datad(rd_ram_rd_addr_1),
	.cin(gnd),
	.combout(\rd_ram_rd_addr[1]~8_combout ),
	.cout());
defparam \rd_ram_rd_addr[1]~8 .lut_mask = 16'h0FF0;
defparam \rd_ram_rd_addr[1]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_rd_addr[2]~9 (
	.dataa(gnd),
	.datab(rd_ram_rd_addr_2),
	.datac(rd_addr_0),
	.datad(rd_ram_rd_addr_1),
	.cin(gnd),
	.combout(\rd_ram_rd_addr[2]~9_combout ),
	.cout());
defparam \rd_ram_rd_addr[2]~9 .lut_mask = 16'hC33C;
defparam \rd_ram_rd_addr[2]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rd_ram_rd_addr[3]~10 (
	.dataa(rd_ram_rd_addr_3),
	.datab(rd_addr_0),
	.datac(rd_ram_rd_addr_1),
	.datad(rd_ram_rd_addr_2),
	.cin(gnd),
	.combout(\rd_ram_rd_addr[3]~10_combout ),
	.cout());
defparam \rd_ram_rd_addr[3]~10 .lut_mask = 16'h6996;
defparam \rd_ram_rd_addr[3]~10 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altsyncram_2 (
	q_b,
	clock1,
	clock0,
	data_a,
	address_a,
	address_b)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	clock1;
input 	clock0;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altsyncram_idh1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clock1(clock1),
	.clock0(clock0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}));

endmodule

module altera_ddr_altsyncram_idh1 (
	q_b,
	clock1,
	clock0,
	data_a,
	address_a,
	address_b)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	clock1;
input 	clock0;
input 	[31:0] data_a;
input 	[3:0] address_a;
input 	[3:0] address_b;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cycloneiii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 4;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 15;
defparam ram_block1a19.port_a_logical_ram_depth = 16;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 4;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 15;
defparam ram_block1a19.port_b_logical_ram_depth = 16;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 4;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 15;
defparam ram_block1a20.port_a_logical_ram_depth = 16;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 4;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 15;
defparam ram_block1a20.port_b_logical_ram_depth = 16;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 4;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 15;
defparam ram_block1a21.port_a_logical_ram_depth = 16;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 4;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 15;
defparam ram_block1a21.port_b_logical_ram_depth = 16;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 4;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 15;
defparam ram_block1a22.port_a_logical_ram_depth = 16;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 4;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 15;
defparam ram_block1a22.port_b_logical_ram_depth = 16;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 4;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 15;
defparam ram_block1a23.port_a_logical_ram_depth = 16;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 4;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 15;
defparam ram_block1a23.port_b_logical_ram_depth = 16;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 4;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 15;
defparam ram_block1a24.port_a_logical_ram_depth = 16;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 4;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 15;
defparam ram_block1a24.port_b_logical_ram_depth = 16;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 4;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 15;
defparam ram_block1a25.port_a_logical_ram_depth = 16;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 4;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 15;
defparam ram_block1a25.port_b_logical_ram_depth = 16;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 4;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 15;
defparam ram_block1a26.port_a_logical_ram_depth = 16;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 4;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 15;
defparam ram_block1a26.port_b_logical_ram_depth = 16;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 4;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 15;
defparam ram_block1a27.port_a_logical_ram_depth = 16;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 4;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 15;
defparam ram_block1a27.port_b_logical_ram_depth = 16;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 4;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 15;
defparam ram_block1a28.port_a_logical_ram_depth = 16;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 4;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 15;
defparam ram_block1a28.port_b_logical_ram_depth = 16;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 4;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 15;
defparam ram_block1a29.port_a_logical_ram_depth = 16;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 4;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 15;
defparam ram_block1a29.port_b_logical_ram_depth = 16;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 4;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 15;
defparam ram_block1a30.port_a_logical_ram_depth = 16;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 4;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 15;
defparam ram_block1a30.port_b_logical_ram_depth = 16;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneiii_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "altera_ddr_controller_phy:altera_ddr_controller_phy_inst|altera_ddr_phy:altera_ddr_phy_inst|altera_ddr_phy_alt_mem_phy:altera_ddr_phy_alt_mem_phy_inst|altera_ddr_phy_alt_mem_phy_read_dp:rdp|altsyncram:full_rate_ram_gen.altsyncram_component|altsyncram_idh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 4;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 15;
defparam ram_block1a31.port_a_logical_ram_depth = 16;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 4;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 15;
defparam ram_block1a31.port_b_logical_ram_depth = 16;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_seq_wrapper (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk_1,
	seq_ac_addr_2,
	seq_ac_addr_3,
	seq_ac_addr_4,
	seq_ac_addr_5,
	dgwb_wdata_24,
	dgwb_wdata_8,
	seq_ac_add_1t_ac_lat_internal,
	ctl_init_success,
	reset_phy_clk_1x_n,
	ctl_init_success1,
	seq_rdv_doing_rd_0,
	seq_rdv_doing_rd_1,
	seq_ac_cs_n_0,
	seq_ac_cke_0,
	seq_ac_addr_0,
	seq_ac_addr_1,
	seq_ac_addr_8,
	seq_ac_addr_10,
	seq_ac_ba_0,
	seq_ac_ba_1,
	seq_ac_ras_n_0,
	seq_ac_cas_n_0,
	seq_ac_we_n_0,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	seq_rdata_valid_lat_dec,
	seq_pll_inc_dec_n,
	seq_pll_start_reconfig,
	seq_mem_clk_disable,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	seq_pll_select_2,
	seq_pll_select_0,
	dgwb_wdata_25,
	dgwb_wdata_9,
	dgwb_wdata_26,
	dgwb_wdata_10,
	dgwb_wdata_27,
	dgwb_wdata_11,
	dgwb_wdata_28,
	dgwb_wdata_12,
	dgwb_wdata_29,
	dgwb_wdata_13,
	dgwb_wdata_30,
	dgwb_wdata_14,
	dgwb_wdata_31,
	dgwb_wdata_15,
	seq_rdata_valid_0,
	phs_shft_busy,
	mimic_done_out,
	seq_mmc_start,
	mimic_value_captured,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	clk_1;
output 	seq_ac_addr_2;
output 	seq_ac_addr_3;
output 	seq_ac_addr_4;
output 	seq_ac_addr_5;
output 	dgwb_wdata_24;
output 	dgwb_wdata_8;
output 	seq_ac_add_1t_ac_lat_internal;
output 	ctl_init_success;
input 	reset_phy_clk_1x_n;
output 	ctl_init_success1;
output 	seq_rdv_doing_rd_0;
output 	seq_rdv_doing_rd_1;
output 	seq_ac_cs_n_0;
output 	seq_ac_cke_0;
output 	seq_ac_addr_0;
output 	seq_ac_addr_1;
output 	seq_ac_addr_8;
output 	seq_ac_addr_10;
output 	seq_ac_ba_0;
output 	seq_ac_ba_1;
output 	seq_ac_ras_n_0;
output 	seq_ac_cas_n_0;
output 	seq_ac_we_n_0;
output 	dgwb_wdp_ovride;
output 	seq_wdp_ovride;
output 	seq_rdata_valid_lat_dec;
output 	seq_pll_inc_dec_n;
output 	seq_pll_start_reconfig;
output 	seq_mem_clk_disable;
output 	wd_lat_0;
output 	wd_lat_1;
output 	wd_lat_4;
output 	wd_lat_3;
output 	wd_lat_2;
output 	seq_pll_select_2;
output 	seq_pll_select_0;
output 	dgwb_wdata_25;
output 	dgwb_wdata_9;
output 	dgwb_wdata_26;
output 	dgwb_wdata_10;
output 	dgwb_wdata_27;
output 	dgwb_wdata_11;
output 	dgwb_wdata_28;
output 	dgwb_wdata_12;
output 	dgwb_wdata_29;
output 	dgwb_wdata_13;
output 	dgwb_wdata_30;
output 	dgwb_wdata_14;
output 	dgwb_wdata_31;
output 	dgwb_wdata_15;
input 	seq_rdata_valid_0;
input 	phs_shft_busy;
input 	mimic_done_out;
output 	seq_mmc_start;
input 	mimic_value_captured;
input 	GND_port;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;



altera_ddr_altera_ddr_phy_alt_mem_phy_seq seq_inst(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk(clk_1),
	.seq_ac_addr_2(seq_ac_addr_2),
	.seq_ac_addr_3(seq_ac_addr_3),
	.seq_ac_addr_4(seq_ac_addr_4),
	.seq_ac_addr_5(seq_ac_addr_5),
	.dgwb_wdata_24(dgwb_wdata_24),
	.dgwb_wdata_8(dgwb_wdata_8),
	.seq_ac_add_1t_ac_lat_internal1(seq_ac_add_1t_ac_lat_internal),
	.ctl_init_success1(ctl_init_success),
	.rst_n(reset_phy_clk_1x_n),
	.ctl_init_success2(ctl_init_success1),
	.seq_rdv_doing_rd_0(seq_rdv_doing_rd_0),
	.seq_rdv_doing_rd_1(seq_rdv_doing_rd_1),
	.seq_ac_cs_n_0(seq_ac_cs_n_0),
	.seq_ac_cke_0(seq_ac_cke_0),
	.seq_ac_addr_0(seq_ac_addr_0),
	.seq_ac_addr_1(seq_ac_addr_1),
	.seq_ac_addr_8(seq_ac_addr_8),
	.seq_ac_addr_10(seq_ac_addr_10),
	.seq_ac_ba_0(seq_ac_ba_0),
	.seq_ac_ba_1(seq_ac_ba_1),
	.seq_ac_ras_n_0(seq_ac_ras_n_0),
	.seq_ac_cas_n_0(seq_ac_cas_n_0),
	.seq_ac_we_n_0(seq_ac_we_n_0),
	.dgwb_wdp_ovride(dgwb_wdp_ovride),
	.seq_wdp_ovride(seq_wdp_ovride),
	.seq_rdata_valid_lat_dec1(seq_rdata_valid_lat_dec),
	.seq_pll_inc_dec_n1(seq_pll_inc_dec_n),
	.seq_pll_start_reconfig1(seq_pll_start_reconfig),
	.seq_mem_clk_disable1(seq_mem_clk_disable),
	.wd_lat_0(wd_lat_0),
	.wd_lat_1(wd_lat_1),
	.wd_lat_4(wd_lat_4),
	.wd_lat_3(wd_lat_3),
	.wd_lat_2(wd_lat_2),
	.seq_pll_select_2(seq_pll_select_2),
	.seq_pll_select_0(seq_pll_select_0),
	.dgwb_wdata_25(dgwb_wdata_25),
	.dgwb_wdata_9(dgwb_wdata_9),
	.dgwb_wdata_26(dgwb_wdata_26),
	.dgwb_wdata_10(dgwb_wdata_10),
	.dgwb_wdata_27(dgwb_wdata_27),
	.dgwb_wdata_11(dgwb_wdata_11),
	.dgwb_wdata_28(dgwb_wdata_28),
	.dgwb_wdata_12(dgwb_wdata_12),
	.dgwb_wdata_29(dgwb_wdata_29),
	.dgwb_wdata_13(dgwb_wdata_13),
	.dgwb_wdata_30(dgwb_wdata_30),
	.dgwb_wdata_14(dgwb_wdata_14),
	.dgwb_wdata_31(dgwb_wdata_31),
	.dgwb_wdata_15(dgwb_wdata_15),
	.rdata_valid({seq_rdata_valid_0}),
	.seq_pll_phs_shift_busy(phs_shft_busy),
	.mmc_seq_done(mimic_done_out),
	.seq_mmc_start(seq_mmc_start),
	.mimic_value_captured(mimic_value_captured),
	.GND_port(GND_port));

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_seq (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk,
	seq_ac_addr_2,
	seq_ac_addr_3,
	seq_ac_addr_4,
	seq_ac_addr_5,
	dgwb_wdata_24,
	dgwb_wdata_8,
	seq_ac_add_1t_ac_lat_internal1,
	ctl_init_success1,
	rst_n,
	ctl_init_success2,
	seq_rdv_doing_rd_0,
	seq_rdv_doing_rd_1,
	seq_ac_cs_n_0,
	seq_ac_cke_0,
	seq_ac_addr_0,
	seq_ac_addr_1,
	seq_ac_addr_8,
	seq_ac_addr_10,
	seq_ac_ba_0,
	seq_ac_ba_1,
	seq_ac_ras_n_0,
	seq_ac_cas_n_0,
	seq_ac_we_n_0,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	seq_rdata_valid_lat_dec1,
	seq_pll_inc_dec_n1,
	seq_pll_start_reconfig1,
	seq_mem_clk_disable1,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	seq_pll_select_2,
	seq_pll_select_0,
	dgwb_wdata_25,
	dgwb_wdata_9,
	dgwb_wdata_26,
	dgwb_wdata_10,
	dgwb_wdata_27,
	dgwb_wdata_11,
	dgwb_wdata_28,
	dgwb_wdata_12,
	dgwb_wdata_29,
	dgwb_wdata_13,
	dgwb_wdata_30,
	dgwb_wdata_14,
	dgwb_wdata_31,
	dgwb_wdata_15,
	rdata_valid,
	seq_pll_phs_shift_busy,
	mmc_seq_done,
	seq_mmc_start,
	mimic_value_captured,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	clk;
output 	seq_ac_addr_2;
output 	seq_ac_addr_3;
output 	seq_ac_addr_4;
output 	seq_ac_addr_5;
output 	dgwb_wdata_24;
output 	dgwb_wdata_8;
output 	seq_ac_add_1t_ac_lat_internal1;
output 	ctl_init_success1;
input 	rst_n;
output 	ctl_init_success2;
output 	seq_rdv_doing_rd_0;
output 	seq_rdv_doing_rd_1;
output 	seq_ac_cs_n_0;
output 	seq_ac_cke_0;
output 	seq_ac_addr_0;
output 	seq_ac_addr_1;
output 	seq_ac_addr_8;
output 	seq_ac_addr_10;
output 	seq_ac_ba_0;
output 	seq_ac_ba_1;
output 	seq_ac_ras_n_0;
output 	seq_ac_cas_n_0;
output 	seq_ac_we_n_0;
output 	dgwb_wdp_ovride;
output 	seq_wdp_ovride;
output 	seq_rdata_valid_lat_dec1;
output 	seq_pll_inc_dec_n1;
output 	seq_pll_start_reconfig1;
output 	seq_mem_clk_disable1;
output 	wd_lat_0;
output 	wd_lat_1;
output 	wd_lat_4;
output 	wd_lat_3;
output 	wd_lat_2;
output 	seq_pll_select_2;
output 	seq_pll_select_0;
output 	dgwb_wdata_25;
output 	dgwb_wdata_9;
output 	dgwb_wdata_26;
output 	dgwb_wdata_10;
output 	dgwb_wdata_27;
output 	dgwb_wdata_11;
output 	dgwb_wdata_28;
output 	dgwb_wdata_12;
output 	dgwb_wdata_29;
output 	dgwb_wdata_13;
output 	dgwb_wdata_30;
output 	dgwb_wdata_14;
output 	dgwb_wdata_31;
output 	dgwb_wdata_15;
input 	[0:0] rdata_valid;
input 	seq_pll_phs_shift_busy;
input 	mmc_seq_done;
output 	seq_mmc_start;
input 	mimic_value_captured;
input 	GND_port;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \admin|addr_cmd[0].cke[0]~q ;
wire \dgwb|sig_addr_cmd[0].addr[2]~q ;
wire \dgwb|sig_addr_cmd[0].addr[3]~q ;
wire \dgwb|sig_addr_cmd[0].addr[4]~q ;
wire \dgwb|sig_addr_cmd[0].addr[5]~q ;
wire \dgwb|sig_addr_cmd[0].cas_n~q ;
wire \pll_ctrl:pll_set_delay[2]~q ;
wire \pll_ctrl:pll_set_delay[1]~q ;
wire \pll_ctrl:pll_set_delay[3]~q ;
wire \pll_ctrl:static_rst_offset[4]~q ;
wire \pll_ctrl:pll_set_delay[1]~3_combout ;
wire \pll_ctrl:pll_set_delay[2]~1_combout ;
wire \pll_ctrl:pll_set_delay[3]~1_combout ;
wire \pll_ctrl:static_rst_offset[4]~1_combout ;
wire \dgrb|sig_doing_rd[0]~q ;
wire \dgrb|sig_doing_rd[1]~q ;
wire \admin|ac_access_gnt~q ;
wire \dgrb|dgrb_ac_access_req~q ;
wire \admin|addr_cmd[0].cs_n[0]~q ;
wire \dgrb|sig_addr_cmd[0].cs_n[0]~q ;
wire \dgwb|dgwb_ac_access_req~q ;
wire \dgwb|sig_addr_cmd[0].cs_n[0]~q ;
wire \admin|addr_cmd[0].addr[0]~q ;
wire \admin|addr_cmd[0].addr[1]~q ;
wire \dgrb|sig_addr_cmd[0].addr[2]~q ;
wire \dgrb|sig_addr_cmd[0].addr[3]~q ;
wire \admin|addr_cmd[0].addr[4]~q ;
wire \dgrb|sig_addr_cmd[0].addr[4]~q ;
wire \dgrb|sig_addr_cmd[0].addr[5]~q ;
wire \admin|addr_cmd[0].addr[8]~q ;
wire \admin|addr_cmd[0].addr[10]~q ;
wire \admin|addr_cmd[0].ba[0]~q ;
wire \admin|addr_cmd[0].ba[1]~q ;
wire \admin|addr_cmd[0].ras_n~q ;
wire \admin|addr_cmd[0].cas_n~q ;
wire \dgrb|sig_addr_cmd[0].cas_n~q ;
wire \admin|addr_cmd[0].we_n~q ;
wire \dgb_ac_access_gnt_r~q ;
wire \dgrb|seq_rdata_valid_lat_dec~q ;
wire \pll_ctrl:pll_set_delay[0]~q ;
wire \Equal1~0_combout ;
wire \pll_ctrl:static_rst_offset[0]~q ;
wire \dgrb|seq_pll_inc_dec_n~q ;
wire \ctrl|state.s_init_dram~q ;
wire \ctrl|WideOr34~8_combout ;
wire \dgrb|seq_pll_start_reconfig~q ;
wire \admin|admin_ctrl.command_done~q ;
wire \dgwb|dgwb_ctrl.command_done~q ;
wire \ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ;
wire \ctrl|Selector1~0_combout ;
wire \ctrl|curr_cmd.cmd_write_btp~q ;
wire \ctrl|curr_cmd.cmd_write_mtp~q ;
wire \ctrl|curr_cmd.cmd_was~q ;
wire \ctrl|WideOr0~0_combout ;
wire \dgrb|dgrb_ctrl.command_done~q ;
wire \ctrl|curr_cmd.cmd_idle~q ;
wire \ctrl|WideOr1~combout ;
wire \ctrl|last_state.s_rdv~q ;
wire \ctrl|last_state.s_read_mtp~q ;
wire \ctrl|last_state.s_rrp_seek~q ;
wire \ctrl|last_state.s_adv_rd_lat~q ;
wire \ctrl|last_state.s_rrp_sweep~q ;
wire \ctrl|last_state.s_adv_wr_lat~q ;
wire \ctrl|last_state.s_rrp_reset~q ;
wire \pll_ctrl:pll_set_delay[0]~0_combout ;
wire \pll_ctrl:static_rst_offset[0]~0_combout ;
wire \dgrb|seq_pll_select[2]~q ;
wire \dgrb|seq_pll_select[0]~q ;
wire \dgb_ac_access_req~0_combout ;
wire \ctrl|Selector58~0_combout ;
wire \ctrl|ctrl_op_rec.command_op.single_bit~0_combout ;
wire \ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ;
wire \ctrl|Selector57~0_combout ;
wire \ctrl|Selector52~0_combout ;
wire \dgrb_phs_shft_busy~q ;
wire \dgrb|dgrb_ctrl.command_result[5]~q ;
wire \dgrb|dgrb_ctrl.command_result[4]~q ;
wire \dgrb|dgrb_ctrl.command_result[3]~q ;
wire \dgrb|dgrb_ctrl.command_result[2]~q ;
wire \dgrb|dgrb_ctrl.command_result[1]~q ;
wire \dgrb|dgrb_ctrl.command_result[0]~q ;
wire \dgrb_phs_shft_busy~2_combout ;
wire \process_4~1_combout ;
wire \seq_ac_addr[2]~13_combout ;
wire \process_4~0_combout ;
wire \seq_ac_addr[3]~14_combout ;
wire \seq_ac_addr[4]~15_combout ;
wire \seq_ac_addr[5]~16_combout ;
wire \seq_ac_cs_n~1_combout ;
wire \seq_ac_cs_n~2_combout ;
wire \v_seq_ac_mux~45_combout ;
wire \seq_ac_cke~1_combout ;
wire \seq_ac_addr~17_combout ;
wire \seq_ac_addr~18_combout ;
wire \seq_ac_addr~19_combout ;
wire \seq_ac_addr~20_combout ;
wire \seq_ac_ba~2_combout ;
wire \seq_ac_ba~3_combout ;
wire \seq_ac_ras_n~1_combout ;
wire \seq_ac_cas_n~3_combout ;
wire \seq_ac_we_n~1_combout ;
wire \seq_ac_cas_n~4_combout ;
wire \seq_ac_we_n~2_combout ;
wire \pll_ctrl:static_rst_offset[1]~2_cout ;
wire \pll_ctrl:static_rst_offset[1]~3_combout ;
wire \pll_ctrl:static_rst_offset[1]~4 ;
wire \pll_ctrl:static_rst_offset[2]~2 ;
wire \pll_ctrl:static_rst_offset[3]~2 ;
wire \pll_ctrl:static_rst_offset[4]~2 ;
wire \pll_ctrl:static_rst_offset[5]~1_combout ;
wire \pll_ctrl:static_rst_offset[5]~q ;
wire \pll_ctrl:static_rst_offset[5]~2 ;
wire \pll_ctrl:static_rst_offset[6]~1_combout ;
wire \pll_ctrl:static_rst_offset[6]~q ;
wire \pll_ctrl:static_rst_offset[6]~2 ;
wire \pll_ctrl:static_rst_offset[7]~3_combout ;
wire \pll_ctrl:static_rst_offset[7]~q ;
wire \Equal0~1_combout ;
wire \seq_pll_phs_shift_busy_r~q ;
wire \seq_pll_phs_shift_busy_ccd~q ;
wire \pll_ctrl:static_rst_offset[7]~1_combout ;
wire \pll_ctrl:static_rst_offset[7]~2_combout ;
wire \pll_ctrl:static_rst_offset[1]~q ;
wire \pll_ctrl:static_rst_offset[2]~1_combout ;
wire \pll_ctrl:static_rst_offset[2]~q ;
wire \pll_ctrl:static_rst_offset[3]~1_combout ;
wire \pll_ctrl:static_rst_offset[3]~q ;
wire \Equal0~0_combout ;
wire \process_13~0_combout ;
wire \seq_pll_inc_dec_n~2_combout ;
wire \pll_ctrl:pll_set_delay[1]~2_cout ;
wire \pll_ctrl:pll_set_delay[1]~4 ;
wire \pll_ctrl:pll_set_delay[2]~2 ;
wire \pll_ctrl:pll_set_delay[3]~2 ;
wire \pll_ctrl:pll_set_delay[4]~2 ;
wire \pll_ctrl:pll_set_delay[5]~1_combout ;
wire \pll_ctrl:pll_set_delay[5]~q ;
wire \pll_ctrl:pll_set_delay[5]~2 ;
wire \pll_ctrl:pll_set_delay[6]~1_combout ;
wire \pll_ctrl:pll_set_delay[6]~q ;
wire \pll_ctrl:pll_set_delay[4]~1_combout ;
wire \pll_ctrl:pll_set_delay[4]~q ;
wire \Equal1~1_combout ;
wire \seq_pll_start_reconfig~3_combout ;
wire \pll_ctrl:phs_shft_busy_1r~0_combout ;
wire \pll_ctrl:phs_shft_busy_1r~q ;
wire \seq_pll_start_reconfig~4_combout ;
wire \ac_mux:ctrl_broadcast_r.command_req~q ;
wire \ac_mux:ctrl_broadcast_r.command.cmd_init_dram~q ;
wire \seq_mem_clk_disable~2_combout ;
wire \seq_pll_select~6_combout ;
wire \seq_pll_select~7_combout ;


altera_ddr_altera_ddr_phy_alt_mem_phy_ctrl ctrl(
	.clk(clk),
	.rst_n(rst_n),
	.ctl_init_success1(ctl_init_success2),
	.states_init_dram(\ctrl|state.s_init_dram~q ),
	.WideOr34(\ctrl|WideOr34~8_combout ),
	.ac_muxctrl_broadcast_rcommandcmd_init_dram(\ac_mux:ctrl_broadcast_r.command.cmd_init_dram~q ),
	.admin_ctrlcommand_done(\admin|admin_ctrl.command_done~q ),
	.dgwb_ctrlcommand_done(\dgwb|dgwb_ctrl.command_done~q ),
	.curr_cmdcmd_prep_customer_mr_setup(\ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ),
	.Selector1(\ctrl|Selector1~0_combout ),
	.curr_cmdcmd_write_btp(\ctrl|curr_cmd.cmd_write_btp~q ),
	.curr_cmdcmd_write_mtp(\ctrl|curr_cmd.cmd_write_mtp~q ),
	.curr_cmdcmd_was(\ctrl|curr_cmd.cmd_was~q ),
	.WideOr0(\ctrl|WideOr0~0_combout ),
	.dgrb_ctrlcommand_done(\dgrb|dgrb_ctrl.command_done~q ),
	.curr_cmdcmd_idle(\ctrl|curr_cmd.cmd_idle~q ),
	.WideOr11(\ctrl|WideOr1~combout ),
	.last_states_rdv(\ctrl|last_state.s_rdv~q ),
	.last_states_read_mtp(\ctrl|last_state.s_read_mtp~q ),
	.last_states_rrp_seek(\ctrl|last_state.s_rrp_seek~q ),
	.last_states_adv_rd_lat(\ctrl|last_state.s_adv_rd_lat~q ),
	.last_states_rrp_sweep(\ctrl|last_state.s_rrp_sweep~q ),
	.last_states_adv_wr_lat(\ctrl|last_state.s_adv_wr_lat~q ),
	.last_states_rrp_reset(\ctrl|last_state.s_rrp_reset~q ),
	.Selector58(\ctrl|Selector58~0_combout ),
	.ctrl_op_reccommand_opsingle_bit(\ctrl|ctrl_op_rec.command_op.single_bit~0_combout ),
	.ctrl_op_reccommand_opmtp_almt(\ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ),
	.Selector57(\ctrl|Selector57~0_combout ),
	.Selector52(\ctrl|Selector52~0_combout ),
	.dgrb_ctrlcommand_result_5(\dgrb|dgrb_ctrl.command_result[5]~q ),
	.dgrb_ctrlcommand_result_4(\dgrb|dgrb_ctrl.command_result[4]~q ),
	.dgrb_ctrlcommand_result_3(\dgrb|dgrb_ctrl.command_result[3]~q ),
	.dgrb_ctrlcommand_result_2(\dgrb|dgrb_ctrl.command_result[2]~q ),
	.dgrb_ctrlcommand_result_1(\dgrb|dgrb_ctrl.command_result[1]~q ),
	.dgrb_ctrlcommand_result_0(\dgrb|dgrb_ctrl.command_result[0]~q ),
	.GND_port(GND_port));

altera_ddr_altera_ddr_phy_alt_mem_phy_admin admin(
	.clk(clk),
	.addr_cmd0cke0(\admin|addr_cmd[0].cke[0]~q ),
	.rst_n(rst_n),
	.ctl_init_success(ctl_init_success2),
	.ac_access_gnt1(\admin|ac_access_gnt~q ),
	.dgrb_ac_access_req(\dgrb|dgrb_ac_access_req~q ),
	.addr_cmd0cs_n0(\admin|addr_cmd[0].cs_n[0]~q ),
	.dgwb_ac_access_req(\dgwb|dgwb_ac_access_req~q ),
	.addr_cmd0addr0(\admin|addr_cmd[0].addr[0]~q ),
	.addr_cmd0addr1(\admin|addr_cmd[0].addr[1]~q ),
	.addr_cmd0addr4(\admin|addr_cmd[0].addr[4]~q ),
	.addr_cmd0addr8(\admin|addr_cmd[0].addr[8]~q ),
	.addr_cmd0addr10(\admin|addr_cmd[0].addr[10]~q ),
	.addr_cmd0ba0(\admin|addr_cmd[0].ba[0]~q ),
	.addr_cmd0ba1(\admin|addr_cmd[0].ba[1]~q ),
	.addr_cmd0ras_n(\admin|addr_cmd[0].ras_n~q ),
	.addr_cmd0cas_n(\admin|addr_cmd[0].cas_n~q ),
	.addr_cmd0we_n(\admin|addr_cmd[0].we_n~q ),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.ac_muxctrl_broadcast_rcommandcmd_init_dram(\ac_mux:ctrl_broadcast_r.command.cmd_init_dram~q ),
	.admin_ctrlcommand_done(\admin|admin_ctrl.command_done~q ),
	.curr_cmdcmd_prep_customer_mr_setup(\ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ),
	.Selector1(\ctrl|Selector1~0_combout ),
	.dgb_ac_access_req(\dgb_ac_access_req~0_combout ),
	.GND_port(GND_port));

altera_ddr_altera_ddr_phy_alt_mem_phy_dgrb dgrb(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_24(q_b_24),
	.q_b_25(q_b_25),
	.q_b_26(q_b_26),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.clk(clk),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal1),
	.rst_n(rst_n),
	.sig_doing_rd_0(\dgrb|sig_doing_rd[0]~q ),
	.sig_doing_rd_1(\dgrb|sig_doing_rd[1]~q ),
	.dgrb_ac_access_req1(\dgrb|dgrb_ac_access_req~q ),
	.sig_addr_cmd0cs_n0(\dgrb|sig_addr_cmd[0].cs_n[0]~q ),
	.sig_addr_cmd0addr2(\dgrb|sig_addr_cmd[0].addr[2]~q ),
	.sig_addr_cmd0addr3(\dgrb|sig_addr_cmd[0].addr[3]~q ),
	.sig_addr_cmd0addr4(\dgrb|sig_addr_cmd[0].addr[4]~q ),
	.sig_addr_cmd0addr5(\dgrb|sig_addr_cmd[0].addr[5]~q ),
	.sig_addr_cmd0cas_n(\dgrb|sig_addr_cmd[0].cas_n~q ),
	.wd_lat_0(wd_lat_0),
	.wd_lat_1(wd_lat_1),
	.wd_lat_4(wd_lat_4),
	.wd_lat_3(wd_lat_3),
	.wd_lat_2(wd_lat_2),
	.dgb_ac_access_gnt_r(\dgb_ac_access_gnt_r~q ),
	.seq_rdata_valid_lat_dec1(\dgrb|seq_rdata_valid_lat_dec~q ),
	.seq_pll_inc_dec_n1(\dgrb|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig1(\dgrb|seq_pll_start_reconfig~q ),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.dgrb_ctrlcommand_done(\dgrb|dgrb_ctrl.command_done~q ),
	.curr_cmdcmd_idle(\ctrl|curr_cmd.cmd_idle~q ),
	.WideOr1(\ctrl|WideOr1~combout ),
	.last_states_rdv(\ctrl|last_state.s_rdv~q ),
	.last_states_read_mtp(\ctrl|last_state.s_read_mtp~q ),
	.last_states_rrp_seek(\ctrl|last_state.s_rrp_seek~q ),
	.last_states_adv_rd_lat(\ctrl|last_state.s_adv_rd_lat~q ),
	.last_states_rrp_sweep(\ctrl|last_state.s_rrp_sweep~q ),
	.last_states_adv_wr_lat(\ctrl|last_state.s_adv_wr_lat~q ),
	.last_states_rrp_reset(\ctrl|last_state.s_rrp_reset~q ),
	.rdata_valid({rdata_valid[0]}),
	.seq_pll_select_2(\dgrb|seq_pll_select[2]~q ),
	.seq_pll_select_0(\dgrb|seq_pll_select[0]~q ),
	.\ctrl_dgrb.command_op.single_bit (\ctrl|ctrl_op_rec.command_op.single_bit~0_combout ),
	.\ctrl_dgrb.command_op.mtp_almt (\ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ),
	.Selector57(\ctrl|Selector57~0_combout ),
	.Selector52(\ctrl|Selector52~0_combout ),
	.phs_shft_busy(\dgrb_phs_shft_busy~q ),
	.dgrb_ctrlcommand_result_5(\dgrb|dgrb_ctrl.command_result[5]~q ),
	.dgrb_ctrlcommand_result_4(\dgrb|dgrb_ctrl.command_result[4]~q ),
	.dgrb_ctrlcommand_result_3(\dgrb|dgrb_ctrl.command_result[3]~q ),
	.dgrb_ctrlcommand_result_2(\dgrb|dgrb_ctrl.command_result[2]~q ),
	.dgrb_ctrlcommand_result_1(\dgrb|dgrb_ctrl.command_result[1]~q ),
	.dgrb_ctrlcommand_result_0(\dgrb|dgrb_ctrl.command_result[0]~q ),
	.mmc_seq_done(mmc_seq_done),
	.seq_mmc_start1(seq_mmc_start),
	.mimic_value_captured(mimic_value_captured),
	.GND_port(GND_port));

altera_ddr_altera_ddr_phy_alt_mem_phy_dgwb dgwb(
	.clk(clk),
	.sig_addr_cmd0addr2(\dgwb|sig_addr_cmd[0].addr[2]~q ),
	.sig_addr_cmd0addr3(\dgwb|sig_addr_cmd[0].addr[3]~q ),
	.sig_addr_cmd0addr4(\dgwb|sig_addr_cmd[0].addr[4]~q ),
	.sig_addr_cmd0addr5(\dgwb|sig_addr_cmd[0].addr[5]~q ),
	.sig_addr_cmd0cas_n(\dgwb|sig_addr_cmd[0].cas_n~q ),
	.dgwb_wdata_24(dgwb_wdata_24),
	.dgwb_wdata_8(dgwb_wdata_8),
	.rst_n(rst_n),
	.dgwb_wdp_ovride1(dgwb_wdp_ovride),
	.dgwb_ac_access_req1(\dgwb|dgwb_ac_access_req~q ),
	.sig_addr_cmd0cs_n0(\dgwb|sig_addr_cmd[0].cs_n[0]~q ),
	.dgb_ac_access_gnt_r(\dgb_ac_access_gnt_r~q ),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.dgwb_ctrlcommand_done(\dgwb|dgwb_ctrl.command_done~q ),
	.curr_cmdcmd_write_btp(\ctrl|curr_cmd.cmd_write_btp~q ),
	.curr_cmdcmd_write_mtp(\ctrl|curr_cmd.cmd_write_mtp~q ),
	.curr_cmdcmd_was(\ctrl|curr_cmd.cmd_was~q ),
	.WideOr0(\ctrl|WideOr0~0_combout ),
	.dgwb_wdata_25(dgwb_wdata_25),
	.dgwb_wdata_9(dgwb_wdata_9),
	.dgwb_wdata_26(dgwb_wdata_26),
	.dgwb_wdata_10(dgwb_wdata_10),
	.dgwb_wdata_27(dgwb_wdata_27),
	.dgwb_wdata_11(dgwb_wdata_11),
	.dgwb_wdata_28(dgwb_wdata_28),
	.dgwb_wdata_12(dgwb_wdata_12),
	.dgwb_wdata_29(dgwb_wdata_29),
	.dgwb_wdata_13(dgwb_wdata_13),
	.dgwb_wdata_30(dgwb_wdata_30),
	.dgwb_wdata_14(dgwb_wdata_14),
	.dgwb_wdata_31(dgwb_wdata_31),
	.dgwb_wdata_15(dgwb_wdata_15));

dffeas \pll_ctrl:pll_set_delay[2] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[2]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[2]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[2] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[2] .power_up = "low";

dffeas \pll_ctrl:pll_set_delay[1] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[1]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[1]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[1] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[1] .power_up = "low";

dffeas \pll_ctrl:pll_set_delay[3] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[3]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[3]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[3] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[3] .power_up = "low";

dffeas \pll_ctrl:static_rst_offset[4] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[4]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[4]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[4] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[4] .power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[1]~3 (
	.dataa(\pll_ctrl:pll_set_delay[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:pll_set_delay[1]~2_cout ),
	.combout(\pll_ctrl:pll_set_delay[1]~3_combout ),
	.cout(\pll_ctrl:pll_set_delay[1]~4 ));
defparam \pll_ctrl:pll_set_delay[1]~3 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:pll_set_delay[1]~3 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[2]~1 (
	.dataa(\pll_ctrl:pll_set_delay[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:pll_set_delay[1]~4 ),
	.combout(\pll_ctrl:pll_set_delay[2]~1_combout ),
	.cout(\pll_ctrl:pll_set_delay[2]~2 ));
defparam \pll_ctrl:pll_set_delay[2]~1 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:pll_set_delay[2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[3]~1 (
	.dataa(\pll_ctrl:pll_set_delay[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:pll_set_delay[2]~2 ),
	.combout(\pll_ctrl:pll_set_delay[3]~1_combout ),
	.cout(\pll_ctrl:pll_set_delay[3]~2 ));
defparam \pll_ctrl:pll_set_delay[3]~1 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:pll_set_delay[3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[4]~1 (
	.dataa(\pll_ctrl:static_rst_offset[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[3]~2 ),
	.combout(\pll_ctrl:static_rst_offset[4]~1_combout ),
	.cout(\pll_ctrl:static_rst_offset[4]~2 ));
defparam \pll_ctrl:static_rst_offset[4]~1 .lut_mask = 16'h5AAF;
defparam \pll_ctrl:static_rst_offset[4]~1 .sum_lutc_input = "cin";

dffeas dgb_ac_access_gnt_r(
	.clk(clk),
	.d(\admin|ac_access_gnt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dgb_ac_access_gnt_r~q ),
	.prn(vcc));
defparam dgb_ac_access_gnt_r.is_wysiwyg = "true";
defparam dgb_ac_access_gnt_r.power_up = "low";

dffeas \pll_ctrl:pll_set_delay[0] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_ctrl:pll_set_delay[0]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[0] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[0] .power_up = "low";

cycloneiii_lcell_comb \Equal1~0 (
	.dataa(\pll_ctrl:pll_set_delay[2]~q ),
	.datab(\pll_ctrl:pll_set_delay[0]~q ),
	.datac(\pll_ctrl:pll_set_delay[1]~q ),
	.datad(\pll_ctrl:pll_set_delay[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hBFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

dffeas \pll_ctrl:static_rst_offset[0] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_ctrl:static_rst_offset[0]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[0] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[0] .power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[0]~0 (
	.dataa(\pll_ctrl:pll_set_delay[0]~q ),
	.datab(\Equal1~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pll_ctrl:pll_set_delay[0]~0_combout ),
	.cout());
defparam \pll_ctrl:pll_set_delay[0]~0 .lut_mask = 16'hDDDD;
defparam \pll_ctrl:pll_set_delay[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[0]~0 (
	.dataa(gnd),
	.datab(\pll_ctrl:static_rst_offset[0]~q ),
	.datac(\pll_ctrl:phs_shft_busy_1r~q ),
	.datad(\pll_ctrl:static_rst_offset[7]~1_combout ),
	.cin(gnd),
	.combout(\pll_ctrl:static_rst_offset[0]~0_combout ),
	.cout());
defparam \pll_ctrl:static_rst_offset[0]~0 .lut_mask = 16'hC33C;
defparam \pll_ctrl:static_rst_offset[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgb_ac_access_req~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\dgwb|dgwb_ac_access_req~q ),
	.datad(\dgrb|dgrb_ac_access_req~q ),
	.cin(gnd),
	.combout(\dgb_ac_access_req~0_combout ),
	.cout());
defparam \dgb_ac_access_req~0 .lut_mask = 16'h0FF0;
defparam \dgb_ac_access_req~0 .sum_lutc_input = "datac";

dffeas dgrb_phs_shft_busy(
	.clk(clk),
	.d(\dgrb_phs_shft_busy~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dgrb_phs_shft_busy~q ),
	.prn(vcc));
defparam dgrb_phs_shft_busy.is_wysiwyg = "true";
defparam dgrb_phs_shft_busy.power_up = "low";

cycloneiii_lcell_comb \dgrb_phs_shft_busy~2 (
	.dataa(\seq_pll_phs_shift_busy_ccd~q ),
	.datab(\seq_pll_start_reconfig~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_phs_shft_busy~2_combout ),
	.cout());
defparam \dgrb_phs_shft_busy~2 .lut_mask = 16'hEEEE;
defparam \dgrb_phs_shft_busy~2 .sum_lutc_input = "datac";

dffeas \seq_ac_addr[2] (
	.clk(clk),
	.d(\seq_ac_addr[2]~13_combout ),
	.asdata(\dgwb|sig_addr_cmd[0].addr[2]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!seq_mem_clk_disable1),
	.sload(\process_4~0_combout ),
	.ena(vcc),
	.q(seq_ac_addr_2),
	.prn(vcc));
defparam \seq_ac_addr[2] .is_wysiwyg = "true";
defparam \seq_ac_addr[2] .power_up = "low";

dffeas \seq_ac_addr[3] (
	.clk(clk),
	.d(\seq_ac_addr[3]~14_combout ),
	.asdata(\dgwb|sig_addr_cmd[0].addr[3]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!seq_mem_clk_disable1),
	.sload(\process_4~0_combout ),
	.ena(vcc),
	.q(seq_ac_addr_3),
	.prn(vcc));
defparam \seq_ac_addr[3] .is_wysiwyg = "true";
defparam \seq_ac_addr[3] .power_up = "low";

dffeas \seq_ac_addr[4] (
	.clk(clk),
	.d(\seq_ac_addr[4]~15_combout ),
	.asdata(\dgwb|sig_addr_cmd[0].addr[4]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!seq_mem_clk_disable1),
	.sload(\process_4~0_combout ),
	.ena(vcc),
	.q(seq_ac_addr_4),
	.prn(vcc));
defparam \seq_ac_addr[4] .is_wysiwyg = "true";
defparam \seq_ac_addr[4] .power_up = "low";

dffeas \seq_ac_addr[5] (
	.clk(clk),
	.d(\seq_ac_addr[5]~16_combout ),
	.asdata(\dgwb|sig_addr_cmd[0].addr[5]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!seq_mem_clk_disable1),
	.sload(\process_4~0_combout ),
	.ena(vcc),
	.q(seq_ac_addr_5),
	.prn(vcc));
defparam \seq_ac_addr[5] .is_wysiwyg = "true";
defparam \seq_ac_addr[5] .power_up = "low";

dffeas seq_ac_add_1t_ac_lat_internal(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_add_1t_ac_lat_internal1),
	.prn(vcc));
defparam seq_ac_add_1t_ac_lat_internal.is_wysiwyg = "true";
defparam seq_ac_add_1t_ac_lat_internal.power_up = "low";

dffeas ctl_init_success(
	.clk(clk),
	.d(ctl_init_success2),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_success1),
	.prn(vcc));
defparam ctl_init_success.is_wysiwyg = "true";
defparam ctl_init_success.power_up = "low";

dffeas \seq_rdv_doing_rd[0] (
	.clk(clk),
	.d(\dgrb|sig_doing_rd[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdv_doing_rd_0),
	.prn(vcc));
defparam \seq_rdv_doing_rd[0] .is_wysiwyg = "true";
defparam \seq_rdv_doing_rd[0] .power_up = "low";

dffeas \seq_rdv_doing_rd[1] (
	.clk(clk),
	.d(\dgrb|sig_doing_rd[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdv_doing_rd_1),
	.prn(vcc));
defparam \seq_rdv_doing_rd[1] .is_wysiwyg = "true";
defparam \seq_rdv_doing_rd[1] .power_up = "low";

dffeas \seq_ac_cs_n[0] (
	.clk(clk),
	.d(\seq_ac_cs_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_cs_n_0),
	.prn(vcc));
defparam \seq_ac_cs_n[0] .is_wysiwyg = "true";
defparam \seq_ac_cs_n[0] .power_up = "low";

dffeas \seq_ac_cke[0] (
	.clk(clk),
	.d(\seq_ac_cke~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_cke_0),
	.prn(vcc));
defparam \seq_ac_cke[0] .is_wysiwyg = "true";
defparam \seq_ac_cke[0] .power_up = "low";

dffeas \seq_ac_addr[0] (
	.clk(clk),
	.d(\seq_ac_addr~17_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_0),
	.prn(vcc));
defparam \seq_ac_addr[0] .is_wysiwyg = "true";
defparam \seq_ac_addr[0] .power_up = "low";

dffeas \seq_ac_addr[1] (
	.clk(clk),
	.d(\seq_ac_addr~18_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_1),
	.prn(vcc));
defparam \seq_ac_addr[1] .is_wysiwyg = "true";
defparam \seq_ac_addr[1] .power_up = "low";

dffeas \seq_ac_addr[8] (
	.clk(clk),
	.d(\seq_ac_addr~19_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_8),
	.prn(vcc));
defparam \seq_ac_addr[8] .is_wysiwyg = "true";
defparam \seq_ac_addr[8] .power_up = "low";

dffeas \seq_ac_addr[10] (
	.clk(clk),
	.d(\seq_ac_addr~20_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_10),
	.prn(vcc));
defparam \seq_ac_addr[10] .is_wysiwyg = "true";
defparam \seq_ac_addr[10] .power_up = "low";

dffeas \seq_ac_ba[0] (
	.clk(clk),
	.d(\seq_ac_ba~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_0),
	.prn(vcc));
defparam \seq_ac_ba[0] .is_wysiwyg = "true";
defparam \seq_ac_ba[0] .power_up = "low";

dffeas \seq_ac_ba[1] (
	.clk(clk),
	.d(\seq_ac_ba~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_1),
	.prn(vcc));
defparam \seq_ac_ba[1] .is_wysiwyg = "true";
defparam \seq_ac_ba[1] .power_up = "low";

dffeas \seq_ac_ras_n[0] (
	.clk(clk),
	.d(\seq_ac_ras_n~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ras_n_0),
	.prn(vcc));
defparam \seq_ac_ras_n[0] .is_wysiwyg = "true";
defparam \seq_ac_ras_n[0] .power_up = "low";

dffeas \seq_ac_cas_n[0] (
	.clk(clk),
	.d(\seq_ac_cas_n~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_cas_n_0),
	.prn(vcc));
defparam \seq_ac_cas_n[0] .is_wysiwyg = "true";
defparam \seq_ac_cas_n[0] .power_up = "low";

dffeas \seq_ac_we_n[0] (
	.clk(clk),
	.d(\seq_ac_we_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_we_n_0),
	.prn(vcc));
defparam \seq_ac_we_n[0] .is_wysiwyg = "true";
defparam \seq_ac_we_n[0] .power_up = "low";

cycloneiii_lcell_comb \seq_wdp_ovride~2 (
	.dataa(dgwb_wdp_ovride),
	.datab(gnd),
	.datac(gnd),
	.datad(ctl_init_success2),
	.cin(gnd),
	.combout(seq_wdp_ovride),
	.cout());
defparam \seq_wdp_ovride~2 .lut_mask = 16'hAAFF;
defparam \seq_wdp_ovride~2 .sum_lutc_input = "datac";

dffeas seq_rdata_valid_lat_dec(
	.clk(clk),
	.d(\dgrb|seq_rdata_valid_lat_dec~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_lat_dec1),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec.power_up = "low";

dffeas seq_pll_inc_dec_n(
	.clk(clk),
	.d(\seq_pll_inc_dec_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_inc_dec_n1),
	.prn(vcc));
defparam seq_pll_inc_dec_n.is_wysiwyg = "true";
defparam seq_pll_inc_dec_n.power_up = "low";

dffeas seq_pll_start_reconfig(
	.clk(clk),
	.d(\seq_pll_start_reconfig~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_start_reconfig1),
	.prn(vcc));
defparam seq_pll_start_reconfig.is_wysiwyg = "true";
defparam seq_pll_start_reconfig.power_up = "low";

dffeas seq_mem_clk_disable(
	.clk(clk),
	.d(\seq_mem_clk_disable~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_mem_clk_disable1),
	.prn(vcc));
defparam seq_mem_clk_disable.is_wysiwyg = "true";
defparam seq_mem_clk_disable.power_up = "low";

dffeas \seq_pll_select[2] (
	.clk(clk),
	.d(\seq_pll_select~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_2),
	.prn(vcc));
defparam \seq_pll_select[2] .is_wysiwyg = "true";
defparam \seq_pll_select[2] .power_up = "low";

dffeas \seq_pll_select[0] (
	.clk(clk),
	.d(\seq_pll_select~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_0),
	.prn(vcc));
defparam \seq_pll_select[0] .is_wysiwyg = "true";
defparam \seq_pll_select[0] .power_up = "low";

cycloneiii_lcell_comb \process_4~1 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgrb|dgrb_ac_access_req~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_4~1_combout ),
	.cout());
defparam \process_4~1 .lut_mask = 16'hEEEE;
defparam \process_4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr[2]~13 (
	.dataa(\admin|addr_cmd[0].addr[0]~q ),
	.datab(\dgrb|sig_addr_cmd[0].addr[2]~q ),
	.datac(gnd),
	.datad(\process_4~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr[2]~13_combout ),
	.cout());
defparam \seq_ac_addr[2]~13 .lut_mask = 16'hAACC;
defparam \seq_ac_addr[2]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_4~0 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgwb|dgwb_ac_access_req~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_4~0_combout ),
	.cout());
defparam \process_4~0 .lut_mask = 16'hEEEE;
defparam \process_4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr[3]~14 (
	.dataa(\admin|addr_cmd[0].addr[0]~q ),
	.datab(\dgrb|sig_addr_cmd[0].addr[3]~q ),
	.datac(gnd),
	.datad(\process_4~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr[3]~14_combout ),
	.cout());
defparam \seq_ac_addr[3]~14 .lut_mask = 16'hAACC;
defparam \seq_ac_addr[3]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr[4]~15 (
	.dataa(\admin|addr_cmd[0].addr[4]~q ),
	.datab(\dgrb|sig_addr_cmd[0].addr[4]~q ),
	.datac(gnd),
	.datad(\process_4~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr[4]~15_combout ),
	.cout());
defparam \seq_ac_addr[4]~15 .lut_mask = 16'hAACC;
defparam \seq_ac_addr[4]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr[5]~16 (
	.dataa(\admin|addr_cmd[0].addr[4]~q ),
	.datab(\dgrb|sig_addr_cmd[0].addr[5]~q ),
	.datac(gnd),
	.datad(\process_4~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr[5]~16_combout ),
	.cout());
defparam \seq_ac_addr[5]~16 .lut_mask = 16'hAACC;
defparam \seq_ac_addr[5]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_cs_n~1 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgrb|dgrb_ac_access_req~q ),
	.datac(\admin|addr_cmd[0].cs_n[0]~q ),
	.datad(\dgrb|sig_addr_cmd[0].cs_n[0]~q ),
	.cin(gnd),
	.combout(\seq_ac_cs_n~1_combout ),
	.cout());
defparam \seq_ac_cs_n~1 .lut_mask = 16'h6FFF;
defparam \seq_ac_cs_n~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_cs_n~2 (
	.dataa(\seq_ac_cs_n~1_combout ),
	.datab(\process_4~0_combout ),
	.datac(\dgwb|sig_addr_cmd[0].cs_n[0]~q ),
	.datad(seq_mem_clk_disable1),
	.cin(gnd),
	.combout(\seq_ac_cs_n~2_combout ),
	.cout());
defparam \seq_ac_cs_n~2 .lut_mask = 16'hF7D5;
defparam \seq_ac_cs_n~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_seq_ac_mux~45 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgwb|dgwb_ac_access_req~q ),
	.datac(\dgrb|dgrb_ac_access_req~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\v_seq_ac_mux~45_combout ),
	.cout());
defparam \v_seq_ac_mux~45 .lut_mask = 16'hFEFE;
defparam \v_seq_ac_mux~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_cke~1 (
	.dataa(seq_mem_clk_disable1),
	.datab(seq_ac_add_1t_ac_lat_internal1),
	.datac(\admin|addr_cmd[0].cke[0]~q ),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_cke~1_combout ),
	.cout());
defparam \seq_ac_cke~1 .lut_mask = 16'hFAFC;
defparam \seq_ac_cke~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr~17 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].addr[0]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr~17_combout ),
	.cout());
defparam \seq_ac_addr~17 .lut_mask = 16'hEEFF;
defparam \seq_ac_addr~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr~18 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].addr[1]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr~18_combout ),
	.cout());
defparam \seq_ac_addr~18 .lut_mask = 16'hEEFF;
defparam \seq_ac_addr~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr~19 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].addr[8]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr~19_combout ),
	.cout());
defparam \seq_ac_addr~19 .lut_mask = 16'hEEFF;
defparam \seq_ac_addr~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_addr~20 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].addr[10]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_addr~20_combout ),
	.cout());
defparam \seq_ac_addr~20 .lut_mask = 16'hEEFF;
defparam \seq_ac_addr~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_ba~2 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].ba[0]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_ba~2_combout ),
	.cout());
defparam \seq_ac_ba~2 .lut_mask = 16'hEEFF;
defparam \seq_ac_ba~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_ba~3 (
	.dataa(seq_mem_clk_disable1),
	.datab(\admin|addr_cmd[0].ba[1]~q ),
	.datac(gnd),
	.datad(\v_seq_ac_mux~45_combout ),
	.cin(gnd),
	.combout(\seq_ac_ba~3_combout ),
	.cout());
defparam \seq_ac_ba~3 .lut_mask = 16'hEEFF;
defparam \seq_ac_ba~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_ras_n~1 (
	.dataa(\v_seq_ac_mux~45_combout ),
	.datab(gnd),
	.datac(seq_mem_clk_disable1),
	.datad(\admin|addr_cmd[0].ras_n~q ),
	.cin(gnd),
	.combout(\seq_ac_ras_n~1_combout ),
	.cout());
defparam \seq_ac_ras_n~1 .lut_mask = 16'hFFF5;
defparam \seq_ac_ras_n~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_cas_n~3 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgrb|dgrb_ac_access_req~q ),
	.datac(\admin|addr_cmd[0].cas_n~q ),
	.datad(\dgrb|sig_addr_cmd[0].cas_n~q ),
	.cin(gnd),
	.combout(\seq_ac_cas_n~3_combout ),
	.cout());
defparam \seq_ac_cas_n~3 .lut_mask = 16'h6FFF;
defparam \seq_ac_cas_n~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_we_n~1 (
	.dataa(seq_mem_clk_disable1),
	.datab(\dgwb|sig_addr_cmd[0].cas_n~q ),
	.datac(\admin|ac_access_gnt~q ),
	.datad(\dgwb|dgwb_ac_access_req~q ),
	.cin(gnd),
	.combout(\seq_ac_we_n~1_combout ),
	.cout());
defparam \seq_ac_we_n~1 .lut_mask = 16'hEFFF;
defparam \seq_ac_we_n~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_cas_n~4 (
	.dataa(\admin|ac_access_gnt~q ),
	.datab(\dgwb|dgwb_ac_access_req~q ),
	.datac(\seq_ac_cas_n~3_combout ),
	.datad(\seq_ac_we_n~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_cas_n~4_combout ),
	.cout());
defparam \seq_ac_cas_n~4 .lut_mask = 16'hFFEF;
defparam \seq_ac_cas_n~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_ac_we_n~2 (
	.dataa(\process_4~1_combout ),
	.datab(\admin|addr_cmd[0].we_n~q ),
	.datac(\process_4~0_combout ),
	.datad(\seq_ac_we_n~1_combout ),
	.cin(gnd),
	.combout(\seq_ac_we_n~2_combout ),
	.cout());
defparam \seq_ac_we_n~2 .lut_mask = 16'hFFFD;
defparam \seq_ac_we_n~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[1]~2 (
	.dataa(\pll_ctrl:static_rst_offset[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\pll_ctrl:static_rst_offset[1]~2_cout ));
defparam \pll_ctrl:static_rst_offset[1]~2 .lut_mask = 16'h00AA;
defparam \pll_ctrl:static_rst_offset[1]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[1]~3 (
	.dataa(\pll_ctrl:static_rst_offset[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[1]~2_cout ),
	.combout(\pll_ctrl:static_rst_offset[1]~3_combout ),
	.cout(\pll_ctrl:static_rst_offset[1]~4 ));
defparam \pll_ctrl:static_rst_offset[1]~3 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:static_rst_offset[1]~3 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[2]~1 (
	.dataa(\pll_ctrl:static_rst_offset[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[1]~4 ),
	.combout(\pll_ctrl:static_rst_offset[2]~1_combout ),
	.cout(\pll_ctrl:static_rst_offset[2]~2 ));
defparam \pll_ctrl:static_rst_offset[2]~1 .lut_mask = 16'h5AAF;
defparam \pll_ctrl:static_rst_offset[2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[3]~1 (
	.dataa(\pll_ctrl:static_rst_offset[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[2]~2 ),
	.combout(\pll_ctrl:static_rst_offset[3]~1_combout ),
	.cout(\pll_ctrl:static_rst_offset[3]~2 ));
defparam \pll_ctrl:static_rst_offset[3]~1 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:static_rst_offset[3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[5]~1 (
	.dataa(\pll_ctrl:static_rst_offset[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[4]~2 ),
	.combout(\pll_ctrl:static_rst_offset[5]~1_combout ),
	.cout(\pll_ctrl:static_rst_offset[5]~2 ));
defparam \pll_ctrl:static_rst_offset[5]~1 .lut_mask = 16'h5A5F;
defparam \pll_ctrl:static_rst_offset[5]~1 .sum_lutc_input = "cin";

dffeas \pll_ctrl:static_rst_offset[5] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[5]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[5]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[5] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[5] .power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[6]~1 (
	.dataa(\pll_ctrl:static_rst_offset[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:static_rst_offset[5]~2 ),
	.combout(\pll_ctrl:static_rst_offset[6]~1_combout ),
	.cout(\pll_ctrl:static_rst_offset[6]~2 ));
defparam \pll_ctrl:static_rst_offset[6]~1 .lut_mask = 16'h5AAF;
defparam \pll_ctrl:static_rst_offset[6]~1 .sum_lutc_input = "cin";

dffeas \pll_ctrl:static_rst_offset[6] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[6]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[6]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[6] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[6] .power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[7]~3 (
	.dataa(\pll_ctrl:static_rst_offset[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\pll_ctrl:static_rst_offset[6]~2 ),
	.combout(\pll_ctrl:static_rst_offset[7]~3_combout ),
	.cout());
defparam \pll_ctrl:static_rst_offset[7]~3 .lut_mask = 16'h5A5A;
defparam \pll_ctrl:static_rst_offset[7]~3 .sum_lutc_input = "cin";

dffeas \pll_ctrl:static_rst_offset[7] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[7]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[7]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[7] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[7] .power_up = "low";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\pll_ctrl:static_rst_offset[4]~q ),
	.datab(\pll_ctrl:static_rst_offset[5]~q ),
	.datac(\pll_ctrl:static_rst_offset[6]~q ),
	.datad(\pll_ctrl:static_rst_offset[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

dffeas seq_pll_phs_shift_busy_r(
	.clk(clk),
	.d(seq_pll_phs_shift_busy),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_phs_shift_busy_r~q ),
	.prn(vcc));
defparam seq_pll_phs_shift_busy_r.is_wysiwyg = "true";
defparam seq_pll_phs_shift_busy_r.power_up = "low";

dffeas seq_pll_phs_shift_busy_ccd(
	.clk(clk),
	.d(\seq_pll_phs_shift_busy_r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_phs_shift_busy_ccd~q ),
	.prn(vcc));
defparam seq_pll_phs_shift_busy_ccd.is_wysiwyg = "true";
defparam seq_pll_phs_shift_busy_ccd.power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[7]~1 (
	.dataa(\Equal1~1_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\seq_pll_phs_shift_busy_ccd~q ),
	.cin(gnd),
	.combout(\pll_ctrl:static_rst_offset[7]~1_combout ),
	.cout());
defparam \pll_ctrl:static_rst_offset[7]~1 .lut_mask = 16'h7FFF;
defparam \pll_ctrl:static_rst_offset[7]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:static_rst_offset[7]~2 (
	.dataa(\pll_ctrl:phs_shft_busy_1r~q ),
	.datab(\pll_ctrl:static_rst_offset[7]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.cout());
defparam \pll_ctrl:static_rst_offset[7]~2 .lut_mask = 16'hEEEE;
defparam \pll_ctrl:static_rst_offset[7]~2 .sum_lutc_input = "datac";

dffeas \pll_ctrl:static_rst_offset[1] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[1]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[1]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[1] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[1] .power_up = "low";

dffeas \pll_ctrl:static_rst_offset[2] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[2]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[2]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[2] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[2] .power_up = "low";

dffeas \pll_ctrl:static_rst_offset[3] (
	.clk(clk),
	.d(\pll_ctrl:static_rst_offset[3]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_ctrl:static_rst_offset[7]~2_combout ),
	.q(\pll_ctrl:static_rst_offset[3]~q ),
	.prn(vcc));
defparam \pll_ctrl:static_rst_offset[3] .is_wysiwyg = "true";
defparam \pll_ctrl:static_rst_offset[3] .power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\pll_ctrl:static_rst_offset[0]~q ),
	.datab(\pll_ctrl:static_rst_offset[1]~q ),
	.datac(\pll_ctrl:static_rst_offset[2]~q ),
	.datad(\pll_ctrl:static_rst_offset[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_13~0 (
	.dataa(\Equal1~1_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\process_13~0_combout ),
	.cout());
defparam \process_13~0 .lut_mask = 16'h5FFF;
defparam \process_13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_inc_dec_n~2 (
	.dataa(\process_13~0_combout ),
	.datab(\dgrb|seq_pll_inc_dec_n~q ),
	.datac(\ctrl|WideOr34~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_pll_inc_dec_n~2_combout ),
	.cout());
defparam \seq_pll_inc_dec_n~2 .lut_mask = 16'hFEFE;
defparam \seq_pll_inc_dec_n~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[1]~2 (
	.dataa(\pll_ctrl:pll_set_delay[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\pll_ctrl:pll_set_delay[1]~2_cout ));
defparam \pll_ctrl:pll_set_delay[1]~2 .lut_mask = 16'h00AA;
defparam \pll_ctrl:pll_set_delay[1]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[4]~1 (
	.dataa(\pll_ctrl:pll_set_delay[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:pll_set_delay[3]~2 ),
	.combout(\pll_ctrl:pll_set_delay[4]~1_combout ),
	.cout(\pll_ctrl:pll_set_delay[4]~2 ));
defparam \pll_ctrl:pll_set_delay[4]~1 .lut_mask = 16'h5AAF;
defparam \pll_ctrl:pll_set_delay[4]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[5]~1 (
	.dataa(\pll_ctrl:pll_set_delay[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pll_ctrl:pll_set_delay[4]~2 ),
	.combout(\pll_ctrl:pll_set_delay[5]~1_combout ),
	.cout(\pll_ctrl:pll_set_delay[5]~2 ));
defparam \pll_ctrl:pll_set_delay[5]~1 .lut_mask = 16'h5AAF;
defparam \pll_ctrl:pll_set_delay[5]~1 .sum_lutc_input = "cin";

dffeas \pll_ctrl:pll_set_delay[5] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[5]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[5]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[5] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[5] .power_up = "low";

cycloneiii_lcell_comb \pll_ctrl:pll_set_delay[6]~1 (
	.dataa(\pll_ctrl:pll_set_delay[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\pll_ctrl:pll_set_delay[5]~2 ),
	.combout(\pll_ctrl:pll_set_delay[6]~1_combout ),
	.cout());
defparam \pll_ctrl:pll_set_delay[6]~1 .lut_mask = 16'h5A5A;
defparam \pll_ctrl:pll_set_delay[6]~1 .sum_lutc_input = "cin";

dffeas \pll_ctrl:pll_set_delay[6] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[6]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[6]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[6] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[6] .power_up = "low";

dffeas \pll_ctrl:pll_set_delay[4] (
	.clk(clk),
	.d(\pll_ctrl:pll_set_delay[4]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal1~1_combout ),
	.q(\pll_ctrl:pll_set_delay[4]~q ),
	.prn(vcc));
defparam \pll_ctrl:pll_set_delay[4] .is_wysiwyg = "true";
defparam \pll_ctrl:pll_set_delay[4] .power_up = "low";

cycloneiii_lcell_comb \Equal1~1 (
	.dataa(\Equal1~0_combout ),
	.datab(\pll_ctrl:pll_set_delay[5]~q ),
	.datac(\pll_ctrl:pll_set_delay[6]~q ),
	.datad(\pll_ctrl:pll_set_delay[4]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hFF7F;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_start_reconfig~3 (
	.dataa(\ctrl|WideOr34~8_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\seq_pll_start_reconfig~3_combout ),
	.cout());
defparam \seq_pll_start_reconfig~3 .lut_mask = 16'hFFFE;
defparam \seq_pll_start_reconfig~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_ctrl:phs_shft_busy_1r~0 (
	.dataa(\seq_pll_phs_shift_busy_ccd~q ),
	.datab(\pll_ctrl:phs_shft_busy_1r~q ),
	.datac(gnd),
	.datad(\process_13~0_combout ),
	.cin(gnd),
	.combout(\pll_ctrl:phs_shft_busy_1r~0_combout ),
	.cout());
defparam \pll_ctrl:phs_shft_busy_1r~0 .lut_mask = 16'hAACC;
defparam \pll_ctrl:phs_shft_busy_1r~0 .sum_lutc_input = "datac";

dffeas \pll_ctrl:phs_shft_busy_1r (
	.clk(clk),
	.d(\pll_ctrl:phs_shft_busy_1r~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_ctrl:phs_shft_busy_1r~q ),
	.prn(vcc));
defparam \pll_ctrl:phs_shft_busy_1r .is_wysiwyg = "true";
defparam \pll_ctrl:phs_shft_busy_1r .power_up = "low";

cycloneiii_lcell_comb \seq_pll_start_reconfig~4 (
	.dataa(\dgrb|seq_pll_start_reconfig~q ),
	.datab(\seq_pll_start_reconfig~3_combout ),
	.datac(\pll_ctrl:static_rst_offset[7]~1_combout ),
	.datad(\pll_ctrl:phs_shft_busy_1r~q ),
	.cin(gnd),
	.combout(\seq_pll_start_reconfig~4_combout ),
	.cout());
defparam \seq_pll_start_reconfig~4 .lut_mask = 16'hFEFF;
defparam \seq_pll_start_reconfig~4 .sum_lutc_input = "datac";

dffeas \ac_mux:ctrl_broadcast_r.command_req (
	.clk(clk),
	.d(\ctrl|Selector58~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.prn(vcc));
defparam \ac_mux:ctrl_broadcast_r.command_req .is_wysiwyg = "true";
defparam \ac_mux:ctrl_broadcast_r.command_req .power_up = "low";

dffeas \ac_mux:ctrl_broadcast_r.command.cmd_init_dram (
	.clk(clk),
	.d(\ctrl|state.s_init_dram~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:ctrl_broadcast_r.command.cmd_init_dram~q ),
	.prn(vcc));
defparam \ac_mux:ctrl_broadcast_r.command.cmd_init_dram .is_wysiwyg = "true";
defparam \ac_mux:ctrl_broadcast_r.command.cmd_init_dram .power_up = "low";

cycloneiii_lcell_comb \seq_mem_clk_disable~2 (
	.dataa(gnd),
	.datab(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.datac(\ac_mux:ctrl_broadcast_r.command.cmd_init_dram~q ),
	.datad(seq_mem_clk_disable1),
	.cin(gnd),
	.combout(\seq_mem_clk_disable~2_combout ),
	.cout());
defparam \seq_mem_clk_disable~2 .lut_mask = 16'hFFFC;
defparam \seq_mem_clk_disable~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_select~6 (
	.dataa(\process_13~0_combout ),
	.datab(\ctrl|WideOr34~8_combout ),
	.datac(\dgrb|seq_pll_select[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_pll_select~6_combout ),
	.cout());
defparam \seq_pll_select~6 .lut_mask = 16'hFEFE;
defparam \seq_pll_select~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_select~7 (
	.dataa(\process_13~0_combout ),
	.datab(\ctrl|WideOr34~8_combout ),
	.datac(\dgrb|seq_pll_select[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_pll_select~7_combout ),
	.cout());
defparam \seq_pll_select~7 .lut_mask = 16'hFEFE;
defparam \seq_pll_select~7 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_admin (
	clk,
	addr_cmd0cke0,
	rst_n,
	ctl_init_success,
	ac_access_gnt1,
	dgrb_ac_access_req,
	addr_cmd0cs_n0,
	dgwb_ac_access_req,
	addr_cmd0addr0,
	addr_cmd0addr1,
	addr_cmd0addr4,
	addr_cmd0addr8,
	addr_cmd0addr10,
	addr_cmd0ba0,
	addr_cmd0ba1,
	addr_cmd0ras_n,
	addr_cmd0cas_n,
	addr_cmd0we_n,
	ac_muxctrl_broadcast_rcommand_req,
	ac_muxctrl_broadcast_rcommandcmd_init_dram,
	admin_ctrlcommand_done,
	curr_cmdcmd_prep_customer_mr_setup,
	Selector1,
	dgb_ac_access_req,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	addr_cmd0cke0;
input 	rst_n;
input 	ctl_init_success;
output 	ac_access_gnt1;
input 	dgrb_ac_access_req;
output 	addr_cmd0cs_n0;
input 	dgwb_ac_access_req;
output 	addr_cmd0addr0;
output 	addr_cmd0addr1;
output 	addr_cmd0addr4;
output 	addr_cmd0addr8;
output 	addr_cmd0addr10;
output 	addr_cmd0ba0;
output 	addr_cmd0ba1;
output 	addr_cmd0ras_n;
output 	addr_cmd0cas_n;
output 	addr_cmd0we_n;
input 	ac_muxctrl_broadcast_rcommand_req;
input 	ac_muxctrl_broadcast_rcommandcmd_init_dram;
output 	admin_ctrlcommand_done;
input 	curr_cmdcmd_prep_customer_mr_setup;
input 	Selector1;
input 	dgb_ac_access_req;
input 	GND_port;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \Add3~22_combout ;
wire \Add3~24_combout ;
wire \Add3~26_combout ;
wire \Add3~34_combout ;
wire \Add3~36_combout ;
wire \Add3~43 ;
wire \Add3~45 ;
wire \Add3~44_combout ;
wire \Add3~47 ;
wire \Add3~46_combout ;
wire \Add3~49 ;
wire \Add3~48_combout ;
wire \Add3~51 ;
wire \Add3~50_combout ;
wire \Add3~53 ;
wire \Add3~52_combout ;
wire \Add3~55 ;
wire \Add3~54_combout ;
wire \Add3~56_combout ;
wire \refresh_count[1]~q ;
wire \refresh_count[2]~q ;
wire \refresh_count[0]~q ;
wire \refresh_count[3]~q ;
wire \refresh_count[6]~q ;
wire \refresh_count[4]~q ;
wire \refresh_count[5]~q ;
wire \refresh_count[7]~q ;
wire \refresh_count[9]~q ;
wire \refresh_count[8]~q ;
wire \refresh_count[0]~31 ;
wire \refresh_count[0]~30_combout ;
wire \refresh_count[1]~33 ;
wire \refresh_count[1]~32_combout ;
wire \initial_refresh_issued~q ;
wire \refresh_count[2]~37 ;
wire \refresh_count[2]~36_combout ;
wire \refresh_count[3]~39 ;
wire \refresh_count[3]~38_combout ;
wire \refresh_count[4]~41 ;
wire \refresh_count[4]~40_combout ;
wire \refresh_count[5]~43 ;
wire \refresh_count[5]~42_combout ;
wire \refresh_count[6]~45 ;
wire \refresh_count[6]~44_combout ;
wire \refresh_count[7]~47 ;
wire \refresh_count[7]~46_combout ;
wire \refresh_count[8]~49 ;
wire \refresh_count[8]~48_combout ;
wire \refresh_count[9]~50_combout ;
wire \Selector302~2_combout ;
wire \Add3~20_combout ;
wire \addr_cmd~513_combout ;
wire \Selector269~3_combout ;
wire \Selector3~0_combout ;
wire \Selector269~4_combout ;
wire \Selector269~5_combout ;
wire \Selector269~7_combout ;
wire \Selector269~8_combout ;
wire \addr_cmd~539_combout ;
wire \addr_cmd~541_combout ;
wire \addr_cmd~542_combout ;
wire \Selector270~1_combout ;
wire \Selector270~2_combout ;
wire \Selector270~3_combout ;
wire \Selector270~4_combout ;
wire \Selector270~5_combout ;
wire \Selector8~0_combout ;
wire \Selector228~0_combout ;
wire \stage_counter[17]~119_combout ;
wire \Selector217~0_combout ;
wire \Selector217~1_combout ;
wire \Selector4~0_combout ;
wire \state~167_combout ;
wire \state~169_combout ;
wire \state~170_combout ;
wire \state~171_combout ;
wire \state~176_combout ;
wire \Selector2~0_combout ;
wire \stage_counter[15]~q ;
wire \stage_counter[14]~q ;
wire \stage_counter[13]~q ;
wire \stage_counter[12]~q ;
wire \stage_counter_zero~1_combout ;
wire \stage_counter[17]~q ;
wire \stage_counter[16]~q ;
wire \stage_counter_zero~2_combout ;
wire \stage_counter[11]~q ;
wire \stage_counter[7]~q ;
wire \Selector221~0_combout ;
wire \Selector3~2_combout ;
wire \Selector249~0_combout ;
wire \finished_state~2_combout ;
wire \stage_counter[0]~q ;
wire \stage_counter[17]~120_combout ;
wire \WideOr26~1_combout ;
wire \stage_counter[17]~122_combout ;
wire \WideNor1~0_combout ;
wire \Add3~58_combout ;
wire \Add3~59_combout ;
wire \Add3~63_combout ;
wire \Add3~64_combout ;
wire \WideNor1~combout ;
wire \stage_counter[5]~128_combout ;
wire \Selector37~0_combout ;
wire \Selector38~0_combout ;
wire \Add3~68_combout ;
wire \Add3~69_combout ;
wire \Add3~73_combout ;
wire \Add3~74_combout ;
wire \Add3~75_combout ;
wire \Add3~76_combout ;
wire \Add3~77_combout ;
wire \Add3~78_combout ;
wire \Add3~81_combout ;
wire \Add3~82_combout ;
wire \Selector10~1_combout ;
wire \Selector249~1_combout ;
wire \stage_counter~138_combout ;
wire \Selector249~2_combout ;
wire \Selector249~3_combout ;
wire \Selector249~4_combout ;
wire \Selector249~5_combout ;
wire \Selector249~6_combout ;
wire \Selector249~7_combout ;
wire \Selector249~8_combout ;
wire \Selector249~9_combout ;
wire \Add3~86_combout ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \refresh_count[1]~34_combout ;
wire \refresh_count[1]~35_combout ;
wire \initial_refresh_issued~2_combout ;
wire \Selector302~5_combout ;
wire \Add3~87_combout ;
wire \Add3~88_combout ;
wire \Add3~89_combout ;
wire \Add3~90_combout ;
wire \Add3~91_combout ;
wire \Add3~92_combout ;
wire \Add3~93_combout ;
wire \state~172_combout ;
wire \state~168_combout ;
wire \Selector15~0_combout ;
wire \command_started~q ;
wire \admin_req_extended~2_combout ;
wire \admin_req_extended~q ;
wire \process_10~0_combout ;
wire \state~173_combout ;
wire \state~175_combout ;
wire \state.s_reset~q ;
wire \state~177_combout ;
wire \state.s_run_init_seq~q ;
wire \addr_cmd[0].cke[0]~0_combout ;
wire \Selector286~2_combout ;
wire \Selector2~1_combout ;
wire \state.s_program_cal_mrs~q ;
wire \WideOr41~0_combout ;
wire \process_7~0_combout ;
wire \refresh_due~q ;
wire \process_8~4_combout ;
wire \num_stacked_refreshes~13_combout ;
wire \num_stacked_refreshes[0]~q ;
wire \process_8~1_combout ;
wire \num_stacked_refreshes~11_combout ;
wire \num_stacked_refreshes~12_combout ;
wire \num_stacked_refreshes[1]~q ;
wire \Selector3~3_combout ;
wire \Selector3~1_combout ;
wire \Selector3~4_combout ;
wire \state~178_combout ;
wire \state.s_access_precharge~q ;
wire \Selector3~5_combout ;
wire \Selector3~6_combout ;
wire \state.s_idle~q ;
wire \Selector216~0_combout ;
wire \Selector216~1_combout ;
wire \Add3~23 ;
wire \Add3~25 ;
wire \Add3~27 ;
wire \Add3~29 ;
wire \Add3~31 ;
wire \Add3~33 ;
wire \Add3~35 ;
wire \Add3~37 ;
wire \Add3~39 ;
wire \Add3~41 ;
wire \Add3~42_combout ;
wire \Add3~94_combout ;
wire \Selector8~1_combout ;
wire \Selector8~2_combout ;
wire \state.s_access~q ;
wire \state~166_combout ;
wire \ac_state.s_10~5_combout ;
wire \ac_state.s_10~3_combout ;
wire \ac_state.s_10~4_combout ;
wire \ac_state.s_10~q ;
wire \Selector228~1_combout ;
wire \ac_state.s_11~q ;
wire \WideOr38~1_combout ;
wire \WideOr41~1_combout ;
wire \ac_state~90_combout ;
wire \ac_state~91_combout ;
wire \ac_state.s_9~q ;
wire \WideOr26~0_combout ;
wire \finished_state~1_combout ;
wire \Selector217~2_combout ;
wire \Selector286~3_combout ;
wire \Selector217~3_combout ;
wire \ac_state.s_0~q ;
wire \process_10~1_combout ;
wire \Selector7~1_combout ;
wire \Selector10~0_combout ;
wire \state.s_prog_user_mrs~q ;
wire \ac_state~93_combout ;
wire \ac_state~94_combout ;
wire \ac_state.s_7~q ;
wire \Add3~21_combout ;
wire \ac_state~95_combout ;
wire \ac_state.s_6~q ;
wire \ac_state~97_combout ;
wire \ac_state.s_5~q ;
wire \process_12~4_combout ;
wire \ac_state~92_combout ;
wire \ac_state.s_8~q ;
wire \process_12~5_combout ;
wire \process_12~6_combout ;
wire \stage_counter[17]~121_combout ;
wire \stage_counter[17]~118_combout ;
wire \Selector269~6_combout ;
wire \stage_counter[17]~123_combout ;
wire \ac_state.s_1~1_combout ;
wire \ac_state.s_1~q ;
wire \state~174_combout ;
wire \state.s_dummy_wait~q ;
wire \WideOr45~1_combout ;
wire \stage_counter[17]~139_combout ;
wire \stage_counter[17]~124_combout ;
wire \stage_counter[17]~125_combout ;
wire \stage_counter[10]~q ;
wire \Add3~40_combout ;
wire \Add3~95_combout ;
wire \stage_counter[9]~q ;
wire \Add3~38_combout ;
wire \Add3~96_combout ;
wire \stage_counter[8]~q ;
wire \stage_counter_zero~3_combout ;
wire \WideOr26~combout ;
wire \stage_counter[5]~126_combout ;
wire \Add3~61_combout ;
wire \Add3~62_combout ;
wire \Add3~65_combout ;
wire \stage_counter[6]~q ;
wire \stage_counter~127_combout ;
wire \Selector19~0_combout ;
wire \stage_counter[5]~129_combout ;
wire \stage_counter[5]~130_combout ;
wire \stage_counter[5]~131_combout ;
wire \stage_counter[5]~132_combout ;
wire \Selector192~0_combout ;
wire \stage_counter~133_combout ;
wire \stage_counter~134_combout ;
wire \Add3~32_combout ;
wire \Add3~66_combout ;
wire \stage_counter[5]~q ;
wire \stage_counter~135_combout ;
wire \Selector20~0_combout ;
wire \Selector193~0_combout ;
wire \stage_counter~136_combout ;
wire \stage_counter~137_combout ;
wire \Add3~30_combout ;
wire \Add3~67_combout ;
wire \stage_counter[4]~q ;
wire \stage_counter_zero~4_combout ;
wire \Add3~70_combout ;
wire \Add3~28_combout ;
wire \Add3~71_combout ;
wire \Add3~72_combout ;
wire \stage_counter[3]~q ;
wire \Add3~60_combout ;
wire \Add3~79_combout ;
wire \Add3~80_combout ;
wire \stage_counter[2]~q ;
wire \Add3~83_combout ;
wire \Add3~84_combout ;
wire \Add3~85_combout ;
wire \stage_counter[1]~q ;
wire \stage_counter_zero~5_combout ;
wire \stage_counter_zero~6_combout ;
wire \stage_counter_zero~q ;
wire \process_12~2_combout ;
wire \per_cs_init_seen[0]~q ;
wire \mem_init_complete~q ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \state.s_topup_refresh~q ;
wire \Selector5~0_combout ;
wire \state.s_topup_refresh_done~q ;
wire \refresh_done~2_combout ;
wire \refresh_done~q ;
wire \num_stacked_refreshes~9_combout ;
wire \num_stacked_refreshes~10_combout ;
wire \num_stacked_refreshes[2]~q ;
wire \LessThan0~0_combout ;
wire \refreshes_maxed~q ;
wire \Selector7~0_combout ;
wire \Selector7~2_combout ;
wire \Selector7~3_combout ;
wire \state.s_access_act~q ;
wire \WideOr43~0_combout ;
wire \Selector219~7_combout ;
wire \Selector219~6_combout ;
wire \ac_state.s_2~q ;
wire \addr_cmd~507_combout ;
wire \finished_state~3_combout ;
wire \finished_state~4_combout ;
wire \finished_state~q ;
wire \Selector13~0_combout ;
wire \state.s_refresh_done~q ;
wire \Selector12~0_combout ;
wire \Selector12~1_combout ;
wire \state.s_refresh~q ;
wire \WideOr45~combout ;
wire \Selector286~5_combout ;
wire \Selector286~4_combout ;
wire \Selector302~3_combout ;
wire \addr_cmd~508_combout ;
wire \Selector302~4_combout ;
wire \Selector269~1_combout ;
wire \addr_cmd~509_combout ;
wire \addr_cmd~510_combout ;
wire \WideNor0~0_combout ;
wire \addr_cmd~511_combout ;
wire \addr_cmd~512_combout ;
wire \Selector269~2_combout ;
wire \Selector269~0_combout ;
wire \addr_cmd~551_combout ;
wire \addr_cmd~514_combout ;
wire \addr_cmd~515_combout ;
wire \addr_cmd~215_combout ;
wire \addr_cmd~516_combout ;
wire \addr_cmd~517_combout ;
wire \addr_cmd~518_combout ;
wire \addr_cmd~519_combout ;
wire \addr_cmd~520_combout ;
wire \addr_cmd~521_combout ;
wire \addr_cmd~522_combout ;
wire \addr_cmd~523_combout ;
wire \addr_cmd~524_combout ;
wire \addr_cmd~525_combout ;
wire \addr_cmd~526_combout ;
wire \addr_cmd~527_combout ;
wire \ac_state~96_combout ;
wire \ac_state.s_3~q ;
wire \Selector221~1_combout ;
wire \ac_state.s_4~q ;
wire \addr_cmd~528_combout ;
wire \addr_cmd~529_combout ;
wire \addr_cmd~530_combout ;
wire \addr_cmd~531_combout ;
wire \addr_cmd~532_combout ;
wire \addr_cmd~533_combout ;
wire \addr_cmd~534_combout ;
wire \addr_cmd~535_combout ;
wire \addr_cmd~536_combout ;
wire \addr_cmd~537_combout ;
wire \Selector269~9_combout ;
wire \addr_cmd~538_combout ;
wire \WideOr32~0_combout ;
wire \addr_cmd~543_combout ;
wire \addr_cmd~540_combout ;
wire \addr_cmd~544_combout ;
wire \addr_cmd~545_combout ;
wire \addr_cmd~546_combout ;
wire \addr_cmd~547_combout ;
wire \addr_cmd~548_combout ;
wire \addr_cmd~549_combout ;
wire \Selector270~0_combout ;
wire \Selector270~6_combout ;
wire \Selector270~7_combout ;
wire \addr_cmd~550_combout ;
wire \command_done~q ;


cycloneiii_lcell_comb \Add3~22 (
	.dataa(\stage_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add3~22_combout ),
	.cout(\Add3~23 ));
defparam \Add3~22 .lut_mask = 16'h55AA;
defparam \Add3~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~24 (
	.dataa(\stage_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~23 ),
	.combout(\Add3~24_combout ),
	.cout(\Add3~25 ));
defparam \Add3~24 .lut_mask = 16'h5A5F;
defparam \Add3~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~26 (
	.dataa(\stage_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~25 ),
	.combout(\Add3~26_combout ),
	.cout(\Add3~27 ));
defparam \Add3~26 .lut_mask = 16'h5AAF;
defparam \Add3~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~34 (
	.dataa(\stage_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~33 ),
	.combout(\Add3~34_combout ),
	.cout(\Add3~35 ));
defparam \Add3~34 .lut_mask = 16'h5AAF;
defparam \Add3~34 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~36 (
	.dataa(\stage_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~35 ),
	.combout(\Add3~36_combout ),
	.cout(\Add3~37 ));
defparam \Add3~36 .lut_mask = 16'h5A5F;
defparam \Add3~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~42 (
	.dataa(\stage_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~41 ),
	.combout(\Add3~42_combout ),
	.cout(\Add3~43 ));
defparam \Add3~42 .lut_mask = 16'h5AAF;
defparam \Add3~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~44 (
	.dataa(\stage_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~43 ),
	.combout(\Add3~44_combout ),
	.cout(\Add3~45 ));
defparam \Add3~44 .lut_mask = 16'h5A5F;
defparam \Add3~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~46 (
	.dataa(\stage_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~45 ),
	.combout(\Add3~46_combout ),
	.cout(\Add3~47 ));
defparam \Add3~46 .lut_mask = 16'h5AAF;
defparam \Add3~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~48 (
	.dataa(\stage_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~47 ),
	.combout(\Add3~48_combout ),
	.cout(\Add3~49 ));
defparam \Add3~48 .lut_mask = 16'h5A5F;
defparam \Add3~48 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~50 (
	.dataa(\stage_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~49 ),
	.combout(\Add3~50_combout ),
	.cout(\Add3~51 ));
defparam \Add3~50 .lut_mask = 16'h5AAF;
defparam \Add3~50 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~52 (
	.dataa(\stage_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~51 ),
	.combout(\Add3~52_combout ),
	.cout(\Add3~53 ));
defparam \Add3~52 .lut_mask = 16'h5A5F;
defparam \Add3~52 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~54 (
	.dataa(\stage_counter[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~53 ),
	.combout(\Add3~54_combout ),
	.cout(\Add3~55 ));
defparam \Add3~54 .lut_mask = 16'h5AAF;
defparam \Add3~54 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~56 (
	.dataa(\stage_counter[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~55 ),
	.combout(\Add3~56_combout ),
	.cout());
defparam \Add3~56 .lut_mask = 16'h5A5A;
defparam \Add3~56 .sum_lutc_input = "cin";

dffeas \refresh_count[1] (
	.clk(clk),
	.d(\refresh_count[1]~32_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[1]~q ),
	.prn(vcc));
defparam \refresh_count[1] .is_wysiwyg = "true";
defparam \refresh_count[1] .power_up = "low";

dffeas \refresh_count[2] (
	.clk(clk),
	.d(\refresh_count[2]~36_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[2]~q ),
	.prn(vcc));
defparam \refresh_count[2] .is_wysiwyg = "true";
defparam \refresh_count[2] .power_up = "low";

dffeas \refresh_count[0] (
	.clk(clk),
	.d(\refresh_count[0]~30_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[0]~q ),
	.prn(vcc));
defparam \refresh_count[0] .is_wysiwyg = "true";
defparam \refresh_count[0] .power_up = "low";

dffeas \refresh_count[3] (
	.clk(clk),
	.d(\refresh_count[3]~38_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[3]~q ),
	.prn(vcc));
defparam \refresh_count[3] .is_wysiwyg = "true";
defparam \refresh_count[3] .power_up = "low";

dffeas \refresh_count[6] (
	.clk(clk),
	.d(\refresh_count[6]~44_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[6]~q ),
	.prn(vcc));
defparam \refresh_count[6] .is_wysiwyg = "true";
defparam \refresh_count[6] .power_up = "low";

dffeas \refresh_count[4] (
	.clk(clk),
	.d(\refresh_count[4]~40_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[4]~q ),
	.prn(vcc));
defparam \refresh_count[4] .is_wysiwyg = "true";
defparam \refresh_count[4] .power_up = "low";

dffeas \refresh_count[5] (
	.clk(clk),
	.d(\refresh_count[5]~42_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[5]~q ),
	.prn(vcc));
defparam \refresh_count[5] .is_wysiwyg = "true";
defparam \refresh_count[5] .power_up = "low";

dffeas \refresh_count[7] (
	.clk(clk),
	.d(\refresh_count[7]~46_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[7]~q ),
	.prn(vcc));
defparam \refresh_count[7] .is_wysiwyg = "true";
defparam \refresh_count[7] .power_up = "low";

dffeas \refresh_count[9] (
	.clk(clk),
	.d(\refresh_count[9]~50_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[9]~q ),
	.prn(vcc));
defparam \refresh_count[9] .is_wysiwyg = "true";
defparam \refresh_count[9] .power_up = "low";

dffeas \refresh_count[8] (
	.clk(clk),
	.d(\refresh_count[8]~48_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\refresh_count[1]~35_combout ),
	.ena(vcc),
	.q(\refresh_count[8]~q ),
	.prn(vcc));
defparam \refresh_count[8] .is_wysiwyg = "true";
defparam \refresh_count[8] .power_up = "low";

cycloneiii_lcell_comb \refresh_count[0]~30 (
	.dataa(\refresh_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\refresh_count[0]~30_combout ),
	.cout(\refresh_count[0]~31 ));
defparam \refresh_count[0]~30 .lut_mask = 16'h55AA;
defparam \refresh_count[0]~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \refresh_count[1]~32 (
	.dataa(\refresh_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[0]~31 ),
	.combout(\refresh_count[1]~32_combout ),
	.cout(\refresh_count[1]~33 ));
defparam \refresh_count[1]~32 .lut_mask = 16'h5AAF;
defparam \refresh_count[1]~32 .sum_lutc_input = "cin";

dffeas initial_refresh_issued(
	.clk(clk),
	.d(\initial_refresh_issued~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\initial_refresh_issued~q ),
	.prn(vcc));
defparam initial_refresh_issued.is_wysiwyg = "true";
defparam initial_refresh_issued.power_up = "low";

cycloneiii_lcell_comb \refresh_count[2]~36 (
	.dataa(\refresh_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[1]~33 ),
	.combout(\refresh_count[2]~36_combout ),
	.cout(\refresh_count[2]~37 ));
defparam \refresh_count[2]~36 .lut_mask = 16'h5A5F;
defparam \refresh_count[2]~36 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[3]~38 (
	.dataa(\refresh_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[2]~37 ),
	.combout(\refresh_count[3]~38_combout ),
	.cout(\refresh_count[3]~39 ));
defparam \refresh_count[3]~38 .lut_mask = 16'h5A5F;
defparam \refresh_count[3]~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[4]~40 (
	.dataa(\refresh_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[3]~39 ),
	.combout(\refresh_count[4]~40_combout ),
	.cout(\refresh_count[4]~41 ));
defparam \refresh_count[4]~40 .lut_mask = 16'h5AAF;
defparam \refresh_count[4]~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[5]~42 (
	.dataa(\refresh_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[4]~41 ),
	.combout(\refresh_count[5]~42_combout ),
	.cout(\refresh_count[5]~43 ));
defparam \refresh_count[5]~42 .lut_mask = 16'h5A5F;
defparam \refresh_count[5]~42 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[6]~44 (
	.dataa(\refresh_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[5]~43 ),
	.combout(\refresh_count[6]~44_combout ),
	.cout(\refresh_count[6]~45 ));
defparam \refresh_count[6]~44 .lut_mask = 16'h5A5F;
defparam \refresh_count[6]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[7]~46 (
	.dataa(\refresh_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[6]~45 ),
	.combout(\refresh_count[7]~46_combout ),
	.cout(\refresh_count[7]~47 ));
defparam \refresh_count[7]~46 .lut_mask = 16'h5A5F;
defparam \refresh_count[7]~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[8]~48 (
	.dataa(\refresh_count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\refresh_count[7]~47 ),
	.combout(\refresh_count[8]~48_combout ),
	.cout(\refresh_count[8]~49 ));
defparam \refresh_count[8]~48 .lut_mask = 16'h5AAF;
defparam \refresh_count[8]~48 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \refresh_count[9]~50 (
	.dataa(\refresh_count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\refresh_count[8]~49 ),
	.combout(\refresh_count[9]~50_combout ),
	.cout());
defparam \refresh_count[9]~50 .lut_mask = 16'h5A5A;
defparam \refresh_count[9]~50 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Selector302~2 (
	.dataa(\WideOr26~combout ),
	.datab(\ac_state.s_0~q ),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\WideOr32~0_combout ),
	.cin(gnd),
	.combout(\Selector302~2_combout ),
	.cout());
defparam \Selector302~2 .lut_mask = 16'hBFFF;
defparam \Selector302~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~20 (
	.dataa(gnd),
	.datab(\ac_state.s_1~q ),
	.datac(\ac_state.s_3~q ),
	.datad(\ac_state.s_4~q ),
	.cin(gnd),
	.combout(\Add3~20_combout ),
	.cout());
defparam \Add3~20 .lut_mask = 16'h3FFF;
defparam \Add3~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~513 (
	.dataa(\addr_cmd~507_combout ),
	.datab(\ac_state.s_1~q ),
	.datac(\state.s_access_act~q ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\addr_cmd~513_combout ),
	.cout());
defparam \addr_cmd~513 .lut_mask = 16'h8BFF;
defparam \addr_cmd~513 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~3 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(addr_cmd0ras_n),
	.datac(\ac_state.s_0~q ),
	.datad(\ac_state.s_8~q ),
	.cin(gnd),
	.combout(\Selector269~3_combout ),
	.cout());
defparam \Selector269~3 .lut_mask = 16'hFEFF;
defparam \Selector269~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\state.s_access_precharge~q ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'h0FFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~4 (
	.dataa(\Selector3~0_combout ),
	.datab(\WideOr45~combout ),
	.datac(\WideOr26~0_combout ),
	.datad(\Selector269~3_combout ),
	.cin(gnd),
	.combout(\Selector269~4_combout ),
	.cout());
defparam \Selector269~4 .lut_mask = 16'hBBF3;
defparam \Selector269~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~5 (
	.dataa(addr_cmd0ras_n),
	.datab(\ac_state.s_0~q ),
	.datac(\state.s_reset~q ),
	.datad(\Selector270~0_combout ),
	.cin(gnd),
	.combout(\Selector269~5_combout ),
	.cout());
defparam \Selector269~5 .lut_mask = 16'hFFFE;
defparam \Selector269~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~7 (
	.dataa(\Selector269~6_combout ),
	.datab(\ac_state.s_1~q ),
	.datac(\Selector270~0_combout ),
	.datad(\Selector269~5_combout ),
	.cin(gnd),
	.combout(\Selector269~7_combout ),
	.cout());
defparam \Selector269~7 .lut_mask = 16'hDFEF;
defparam \Selector269~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~8 (
	.dataa(\Selector269~3_combout ),
	.datab(\Selector269~4_combout ),
	.datac(\Selector269~5_combout ),
	.datad(\Selector269~7_combout ),
	.cin(gnd),
	.combout(\Selector269~8_combout ),
	.cout());
defparam \Selector269~8 .lut_mask = 16'hEBBE;
defparam \Selector269~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~539 (
	.dataa(\state.s_reset~q ),
	.datab(\state.s_access_act~q ),
	.datac(gnd),
	.datad(\ac_state.s_1~q ),
	.cin(gnd),
	.combout(\addr_cmd~539_combout ),
	.cout());
defparam \addr_cmd~539 .lut_mask = 16'hEEFF;
defparam \addr_cmd~539 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~541 (
	.dataa(\ac_state.s_3~q ),
	.datab(\ac_state.s_2~q ),
	.datac(\ac_state.s_5~q ),
	.datad(\addr_cmd~540_combout ),
	.cin(gnd),
	.combout(\addr_cmd~541_combout ),
	.cout());
defparam \addr_cmd~541 .lut_mask = 16'hFFFE;
defparam \addr_cmd~541 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~542 (
	.dataa(addr_cmd0cas_n),
	.datab(\addr_cmd~539_combout ),
	.datac(\addr_cmd~541_combout ),
	.datad(\stage_counter[17]~118_combout ),
	.cin(gnd),
	.combout(\addr_cmd~542_combout ),
	.cout());
defparam \addr_cmd~542 .lut_mask = 16'hFFFE;
defparam \addr_cmd~542 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~1 (
	.dataa(addr_cmd0we_n),
	.datab(\state.s_reset~q ),
	.datac(\WideOr26~0_combout ),
	.datad(\Selector269~0_combout ),
	.cin(gnd),
	.combout(\Selector270~1_combout ),
	.cout());
defparam \Selector270~1 .lut_mask = 16'hEFFF;
defparam \Selector270~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~2 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(\Selector270~1_combout ),
	.datac(\Add3~20_combout ),
	.datad(\Add3~21_combout ),
	.cin(gnd),
	.combout(\Selector270~2_combout ),
	.cout());
defparam \Selector270~2 .lut_mask = 16'hEFFF;
defparam \Selector270~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~3 (
	.dataa(addr_cmd0we_n),
	.datab(\state.s_reset~q ),
	.datac(\WideOr45~1_combout ),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector270~3_combout ),
	.cout());
defparam \Selector270~3 .lut_mask = 16'hEFFF;
defparam \Selector270~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~4 (
	.dataa(\Selector270~2_combout ),
	.datab(\Selector270~3_combout ),
	.datac(addr_cmd0we_n),
	.datad(\WideOr38~1_combout ),
	.cin(gnd),
	.combout(\Selector270~4_combout ),
	.cout());
defparam \Selector270~4 .lut_mask = 16'hFEFF;
defparam \Selector270~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~5 (
	.dataa(addr_cmd0we_n),
	.datab(\state.s_reset~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\Selector269~6_combout ),
	.cin(gnd),
	.combout(\Selector270~5_combout ),
	.cout());
defparam \Selector270~5 .lut_mask = 16'hEFFF;
defparam \Selector270~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~0 (
	.dataa(\state.s_access_act~q ),
	.datab(\finished_state~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hEEEE;
defparam \Selector8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector228~0 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\ac_state.s_10~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector228~0_combout ),
	.cout());
defparam \Selector228~0 .lut_mask = 16'hEEEE;
defparam \Selector228~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~119 (
	.dataa(\state.s_topup_refresh~q ),
	.datab(\state.s_refresh~q ),
	.datac(\state.s_access_act~q ),
	.datad(\state.s_access_precharge~q ),
	.cin(gnd),
	.combout(\stage_counter[17]~119_combout ),
	.cout());
defparam \stage_counter[17]~119 .lut_mask = 16'hFFFE;
defparam \stage_counter[17]~119 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector217~0 (
	.dataa(\ac_state.s_0~q ),
	.datab(\stage_counter[17]~119_combout ),
	.datac(\ac_state.s_1~q ),
	.datad(\WideOr45~1_combout ),
	.cin(gnd),
	.combout(\Selector217~0_combout ),
	.cout());
defparam \Selector217~0 .lut_mask = 16'hEFFF;
defparam \Selector217~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector217~1 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\ac_state.s_7~q ),
	.datac(\WideOr26~combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector217~1_combout ),
	.cout());
defparam \Selector217~1 .lut_mask = 16'hFEFE;
defparam \Selector217~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\state.s_topup_refresh~q ),
	.datab(\Selector7~1_combout ),
	.datac(\state.s_idle~q ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFEFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~167 (
	.dataa(\mem_init_complete~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\refreshes_maxed~q ),
	.cin(gnd),
	.combout(\state~167_combout ),
	.cout());
defparam \state~167 .lut_mask = 16'hAAFF;
defparam \state~167 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~169 (
	.dataa(\state~167_combout ),
	.datab(\state~168_combout ),
	.datac(\process_10~0_combout ),
	.datad(\process_10~1_combout ),
	.cin(gnd),
	.combout(\state~169_combout ),
	.cout());
defparam \state~169 .lut_mask = 16'hEFFF;
defparam \state~169 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~170 (
	.dataa(dgb_ac_access_req),
	.datab(\state~167_combout ),
	.datac(\admin_req_extended~q ),
	.datad(Selector1),
	.cin(gnd),
	.combout(\state~170_combout ),
	.cout());
defparam \state~170 .lut_mask = 16'hFEFF;
defparam \state~170 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~171 (
	.dataa(\state.s_idle~q ),
	.datab(\finished_state~q ),
	.datac(\state~166_combout ),
	.datad(\state~170_combout ),
	.cin(gnd),
	.combout(\state~171_combout ),
	.cout());
defparam \state~171 .lut_mask = 16'hFFFE;
defparam \state~171 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~176 (
	.dataa(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datab(\admin_req_extended~q ),
	.datac(gnd),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\state~176_combout ),
	.cout());
defparam \state~176 .lut_mask = 16'hEEFF;
defparam \state~176 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~0 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(\process_10~0_combout ),
	.datac(\state~168_combout ),
	.datad(\Selector7~1_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFFFE;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \stage_counter[15] (
	.clk(clk),
	.d(\Add3~87_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[15]~q ),
	.prn(vcc));
defparam \stage_counter[15] .is_wysiwyg = "true";
defparam \stage_counter[15] .power_up = "low";

dffeas \stage_counter[14] (
	.clk(clk),
	.d(\Add3~88_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[14]~q ),
	.prn(vcc));
defparam \stage_counter[14] .is_wysiwyg = "true";
defparam \stage_counter[14] .power_up = "low";

dffeas \stage_counter[13] (
	.clk(clk),
	.d(\Add3~89_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[13]~q ),
	.prn(vcc));
defparam \stage_counter[13] .is_wysiwyg = "true";
defparam \stage_counter[13] .power_up = "low";

dffeas \stage_counter[12] (
	.clk(clk),
	.d(\Add3~90_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[12]~q ),
	.prn(vcc));
defparam \stage_counter[12] .is_wysiwyg = "true";
defparam \stage_counter[12] .power_up = "low";

cycloneiii_lcell_comb \stage_counter_zero~1 (
	.dataa(\stage_counter[15]~q ),
	.datab(\stage_counter[14]~q ),
	.datac(\stage_counter[13]~q ),
	.datad(\stage_counter[12]~q ),
	.cin(gnd),
	.combout(\stage_counter_zero~1_combout ),
	.cout());
defparam \stage_counter_zero~1 .lut_mask = 16'h7FFF;
defparam \stage_counter_zero~1 .sum_lutc_input = "datac";

dffeas \stage_counter[17] (
	.clk(clk),
	.d(\Add3~91_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[17]~q ),
	.prn(vcc));
defparam \stage_counter[17] .is_wysiwyg = "true";
defparam \stage_counter[17] .power_up = "low";

dffeas \stage_counter[16] (
	.clk(clk),
	.d(\Add3~92_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[16]~q ),
	.prn(vcc));
defparam \stage_counter[16] .is_wysiwyg = "true";
defparam \stage_counter[16] .power_up = "low";

cycloneiii_lcell_comb \stage_counter_zero~2 (
	.dataa(\stage_counter_zero~1_combout ),
	.datab(\process_12~2_combout ),
	.datac(\stage_counter[17]~q ),
	.datad(\stage_counter[16]~q ),
	.cin(gnd),
	.combout(\stage_counter_zero~2_combout ),
	.cout());
defparam \stage_counter_zero~2 .lut_mask = 16'hBFFF;
defparam \stage_counter_zero~2 .sum_lutc_input = "datac";

dffeas \stage_counter[11] (
	.clk(clk),
	.d(\Add3~93_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[11]~q ),
	.prn(vcc));
defparam \stage_counter[11] .is_wysiwyg = "true";
defparam \stage_counter[11] .power_up = "low";

dffeas \stage_counter[7] (
	.clk(clk),
	.d(\Add3~63_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[7]~q ),
	.prn(vcc));
defparam \stage_counter[7] .is_wysiwyg = "true";
defparam \stage_counter[7] .power_up = "low";

cycloneiii_lcell_comb \Selector221~0 (
	.dataa(\ac_state.s_1~q ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\ac_state.s_4~q ),
	.datad(\state~166_combout ),
	.cin(gnd),
	.combout(\Selector221~0_combout ),
	.cout());
defparam \Selector221~0 .lut_mask = 16'hFEFF;
defparam \Selector221~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~2 (
	.dataa(\state.s_idle~q ),
	.datab(\Selector8~1_combout ),
	.datac(\Selector3~0_combout ),
	.datad(\state~170_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'hEFFF;
defparam \Selector3~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~0 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\ac_state.s_11~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector249~0_combout ),
	.cout());
defparam \Selector249~0 .lut_mask = 16'hEEEE;
defparam \Selector249~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \finished_state~2 (
	.dataa(\finished_state~1_combout ),
	.datab(\Selector249~0_combout ),
	.datac(\ac_state.s_1~q ),
	.datad(\WideOr45~1_combout ),
	.cin(gnd),
	.combout(\finished_state~2_combout ),
	.cout());
defparam \finished_state~2 .lut_mask = 16'hFEFF;
defparam \finished_state~2 .sum_lutc_input = "datac";

dffeas \stage_counter[0] (
	.clk(clk),
	.d(\Add3~86_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[0]~q ),
	.prn(vcc));
defparam \stage_counter[0] .is_wysiwyg = "true";
defparam \stage_counter[0] .power_up = "low";

cycloneiii_lcell_comb \stage_counter[17]~120 (
	.dataa(\state.s_reset~q ),
	.datab(\state.s_access~q ),
	.datac(\stage_counter_zero~q ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\stage_counter[17]~120_combout ),
	.cout());
defparam \stage_counter[17]~120 .lut_mask = 16'hBFFF;
defparam \stage_counter[17]~120 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr26~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_10~q ),
	.datad(\ac_state.s_11~q ),
	.cin(gnd),
	.combout(\WideOr26~1_combout ),
	.cout());
defparam \WideOr26~1 .lut_mask = 16'h0FFF;
defparam \WideOr26~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~122 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\WideOr26~combout ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(\WideOr26~1_combout ),
	.cin(gnd),
	.combout(\stage_counter[17]~122_combout ),
	.cout());
defparam \stage_counter[17]~122 .lut_mask = 16'hACFF;
defparam \stage_counter[17]~122 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~0 (
	.dataa(\ac_state.s_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_state.s_1~q ),
	.cin(gnd),
	.combout(\WideNor1~0_combout ),
	.cout());
defparam \WideNor1~0 .lut_mask = 16'hAAFF;
defparam \WideNor1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~58 (
	.dataa(\ac_state.s_8~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\Add3~58_combout ),
	.cout());
defparam \Add3~58 .lut_mask = 16'hEFFF;
defparam \Add3~58 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~59 (
	.dataa(\Add3~58_combout ),
	.datab(\Selector228~0_combout ),
	.datac(\Add3~36_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~59_combout ),
	.cout());
defparam \Add3~59 .lut_mask = 16'hFAFC;
defparam \Add3~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~63 (
	.dataa(\Add3~59_combout ),
	.datab(\stage_counter[7]~q ),
	.datac(\Add3~62_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~63_combout ),
	.cout());
defparam \Add3~63 .lut_mask = 16'hFEFE;
defparam \Add3~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~64 (
	.dataa(\ac_state.s_8~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\Add3~34_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~64_combout ),
	.cout());
defparam \Add3~64 .lut_mask = 16'hFAFC;
defparam \Add3~64 .sum_lutc_input = "datac";

cycloneiii_lcell_comb WideNor1(
	.dataa(\ac_state.s_0~q ),
	.datab(gnd),
	.datac(\ac_state.s_1~q ),
	.datad(\ac_state.s_2~q ),
	.cin(gnd),
	.combout(\WideNor1~combout ),
	.cout());
defparam WideNor1.lut_mask = 16'hAFFF;
defparam WideNor1.sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~128 (
	.dataa(\WideOr26~combout ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\WideNor1~combout ),
	.datad(\state.s_dummy_wait~q ),
	.cin(gnd),
	.combout(\stage_counter[5]~128_combout ),
	.cout());
defparam \stage_counter[5]~128 .lut_mask = 16'hB8FF;
defparam \stage_counter[5]~128 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector37~0 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[5]~q ),
	.datac(\WideOr26~1_combout ),
	.datad(\process_12~4_combout ),
	.cin(gnd),
	.combout(\Selector37~0_combout ),
	.cout());
defparam \Selector37~0 .lut_mask = 16'hEFFF;
defparam \Selector37~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector38~0 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[4]~q ),
	.datac(\WideOr26~1_combout ),
	.datad(\process_12~4_combout ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hEFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~68 (
	.dataa(\ac_state.s_1~q ),
	.datab(\process_12~2_combout ),
	.datac(\state.s_access_act~q ),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Add3~68_combout ),
	.cout());
defparam \Add3~68 .lut_mask = 16'hFEFF;
defparam \Add3~68 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~69 (
	.dataa(\Add3~68_combout ),
	.datab(\addr_cmd~520_combout ),
	.datac(\ac_state.s_8~q ),
	.datad(\Add3~20_combout ),
	.cin(gnd),
	.combout(\Add3~69_combout ),
	.cout());
defparam \Add3~69 .lut_mask = 16'hFEFF;
defparam \Add3~69 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~73 (
	.dataa(\addr_cmd~532_combout ),
	.datab(\ac_state.s_3~q ),
	.datac(\ac_state.s_4~q ),
	.datad(\ac_state.s_2~q ),
	.cin(gnd),
	.combout(\Add3~73_combout ),
	.cout());
defparam \Add3~73 .lut_mask = 16'hFFFE;
defparam \Add3~73 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~74 (
	.dataa(gnd),
	.datab(\state.s_reset~q ),
	.datac(\stage_counter_zero~q ),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Add3~74_combout ),
	.cout());
defparam \Add3~74 .lut_mask = 16'h3FFF;
defparam \Add3~74 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~75 (
	.dataa(\Add3~73_combout ),
	.datab(\Add3~74_combout ),
	.datac(\state.s_access_act~q ),
	.datad(\WideOr45~1_combout ),
	.cin(gnd),
	.combout(\Add3~75_combout ),
	.cout());
defparam \Add3~75 .lut_mask = 16'hFEFF;
defparam \Add3~75 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~76 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(\process_12~2_combout ),
	.datac(\Add3~21_combout ),
	.datad(\process_12~4_combout ),
	.cin(gnd),
	.combout(\Add3~76_combout ),
	.cout());
defparam \Add3~76 .lut_mask = 16'hEFFF;
defparam \Add3~76 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~77 (
	.dataa(\Add3~75_combout ),
	.datab(\Add3~76_combout ),
	.datac(\Add3~26_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~77_combout ),
	.cout());
defparam \Add3~77 .lut_mask = 16'hFEFF;
defparam \Add3~77 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~78 (
	.dataa(\Add3~77_combout ),
	.datab(\state.s_run_init_seq~q ),
	.datac(\process_12~6_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~78_combout ),
	.cout());
defparam \Add3~78 .lut_mask = 16'hFFFE;
defparam \Add3~78 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~81 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\ac_state.s_10~q ),
	.datac(\Add3~24_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~81_combout ),
	.cout());
defparam \Add3~81 .lut_mask = 16'hFAFC;
defparam \Add3~81 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~82 (
	.dataa(\Add3~81_combout ),
	.datab(\addr_cmd~520_combout ),
	.datac(\process_12~4_combout ),
	.datad(\refresh_done~2_combout ),
	.cin(gnd),
	.combout(\Add3~82_combout ),
	.cout());
defparam \Add3~82 .lut_mask = 16'hFFEF;
defparam \Add3~82 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~1 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\finished_state~q ),
	.datac(\refreshes_maxed~q ),
	.datad(\process_10~1_combout ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hFFFE;
defparam \Selector10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~1 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[0]~q ),
	.datac(\stage_counter[17]~121_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector249~1_combout ),
	.cout());
defparam \Selector249~1 .lut_mask = 16'hFEFE;
defparam \Selector249~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter~138 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter~138_combout ),
	.cout());
defparam \stage_counter~138 .lut_mask = 16'hEEEE;
defparam \stage_counter~138 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~2 (
	.dataa(\ac_state.s_2~q ),
	.datab(\WideNor1~0_combout ),
	.datac(\stage_counter~138_combout ),
	.datad(\WideOr43~0_combout ),
	.cin(gnd),
	.combout(\Selector249~2_combout ),
	.cout());
defparam \Selector249~2 .lut_mask = 16'hFEFF;
defparam \Selector249~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~3 (
	.dataa(\stage_counter~138_combout ),
	.datab(\WideNor1~combout ),
	.datac(\addr_cmd~507_combout ),
	.datad(\state~166_combout ),
	.cin(gnd),
	.combout(\Selector249~3_combout ),
	.cout());
defparam \Selector249~3 .lut_mask = 16'hBFFF;
defparam \Selector249~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~4 (
	.dataa(\ac_state.s_9~q ),
	.datab(\stage_counter~138_combout ),
	.datac(\WideOr26~1_combout ),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Selector249~4_combout ),
	.cout());
defparam \Selector249~4 .lut_mask = 16'hEFFF;
defparam \Selector249~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~5 (
	.dataa(\Selector249~0_combout ),
	.datab(\Selector249~3_combout ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(\Selector249~4_combout ),
	.cin(gnd),
	.combout(\Selector249~5_combout ),
	.cout());
defparam \Selector249~5 .lut_mask = 16'hFFFE;
defparam \Selector249~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~6 (
	.dataa(\WideOr26~combout ),
	.datab(\stage_counter~138_combout ),
	.datac(\ac_state.s_0~q ),
	.datad(\WideOr32~0_combout ),
	.cin(gnd),
	.combout(\Selector249~6_combout ),
	.cout());
defparam \Selector249~6 .lut_mask = 16'hEFFF;
defparam \Selector249~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~7 (
	.dataa(\Selector249~2_combout ),
	.datab(\Selector249~5_combout ),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\Selector249~6_combout ),
	.cin(gnd),
	.combout(\Selector249~7_combout ),
	.cout());
defparam \Selector249~7 .lut_mask = 16'hFFFE;
defparam \Selector249~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~8 (
	.dataa(\ac_state.s_1~q ),
	.datab(\ac_state.s_0~q ),
	.datac(\stage_counter~138_combout ),
	.datad(\WideOr45~1_combout ),
	.cin(gnd),
	.combout(\Selector249~8_combout ),
	.cout());
defparam \Selector249~8 .lut_mask = 16'hFEFF;
defparam \Selector249~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector249~9 (
	.dataa(\Selector249~7_combout ),
	.datab(\Selector249~8_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\Selector249~9_combout ),
	.cout());
defparam \Selector249~9 .lut_mask = 16'hFFFE;
defparam \Selector249~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~86 (
	.dataa(\Add3~22_combout ),
	.datab(\process_12~2_combout ),
	.datac(\Selector249~1_combout ),
	.datad(\Selector249~9_combout ),
	.cin(gnd),
	.combout(\Add3~86_combout ),
	.cout());
defparam \Add3~86 .lut_mask = 16'hFFB8;
defparam \Add3~86 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\refresh_count[1]~q ),
	.datab(\refresh_count[2]~q ),
	.datac(\refresh_count[0]~q ),
	.datad(\refresh_count[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\refresh_count[6]~q ),
	.datab(\refresh_count[4]~q ),
	.datac(\refresh_count[5]~q ),
	.datad(\refresh_count[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hBFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\refresh_count[9]~q ),
	.datad(\refresh_count[8]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \refresh_count[1]~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\refreshes_maxed~q ),
	.datad(\refresh_done~q ),
	.cin(gnd),
	.combout(\refresh_count[1]~34_combout ),
	.cout());
defparam \refresh_count[1]~34 .lut_mask = 16'h0FFF;
defparam \refresh_count[1]~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \refresh_count[1]~35 (
	.dataa(\refresh_count[1]~34_combout ),
	.datab(\initial_refresh_issued~q ),
	.datac(ctl_init_success),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\refresh_count[1]~35_combout ),
	.cout());
defparam \refresh_count[1]~35 .lut_mask = 16'hFFF7;
defparam \refresh_count[1]~35 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \initial_refresh_issued~2 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_refresh_done~q ),
	.datac(\initial_refresh_issued~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\initial_refresh_issued~2_combout ),
	.cout());
defparam \initial_refresh_issued~2 .lut_mask = 16'hFEFE;
defparam \initial_refresh_issued~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector302~5 (
	.dataa(\ac_state.s_0~q ),
	.datab(\ac_state.s_8~q ),
	.datac(\WideOr26~0_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\Selector302~5_combout ),
	.cout());
defparam \Selector302~5 .lut_mask = 16'hDFFF;
defparam \Selector302~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~87 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~87_combout ),
	.cout());
defparam \Add3~87 .lut_mask = 16'hFEFE;
defparam \Add3~87 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~88 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~50_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~88_combout ),
	.cout());
defparam \Add3~88 .lut_mask = 16'hFEFE;
defparam \Add3~88 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~89 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~89_combout ),
	.cout());
defparam \Add3~89 .lut_mask = 16'hFEFE;
defparam \Add3~89 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~90 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~90_combout ),
	.cout());
defparam \Add3~90 .lut_mask = 16'hFEFE;
defparam \Add3~90 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~91 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~56_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~91_combout ),
	.cout());
defparam \Add3~91 .lut_mask = 16'hFEFE;
defparam \Add3~91 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~92 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~54_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~92_combout ),
	.cout());
defparam \Add3~92 .lut_mask = 16'hFEFE;
defparam \Add3~92 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~93 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~93_combout ),
	.cout());
defparam \Add3~93 .lut_mask = 16'hFEFE;
defparam \Add3~93 .sum_lutc_input = "datac";

dffeas \addr_cmd[0].cke[0] (
	.clk(clk),
	.d(\addr_cmd[0].cke[0]~0_combout ),
	.asdata(\Selector286~4_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_12~2_combout ),
	.ena(vcc),
	.q(addr_cmd0cke0),
	.prn(vcc));
defparam \addr_cmd[0].cke[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].cke[0] .power_up = "low";

dffeas ac_access_gnt(
	.clk(clk),
	.d(\state.s_access~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac_access_gnt1),
	.prn(vcc));
defparam ac_access_gnt.is_wysiwyg = "true";
defparam ac_access_gnt.power_up = "low";

dffeas \addr_cmd[0].cs_n[0] (
	.clk(clk),
	.d(\addr_cmd~511_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0cs_n0),
	.prn(vcc));
defparam \addr_cmd[0].cs_n[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].cs_n[0] .power_up = "low";

dffeas \addr_cmd[0].addr[0] (
	.clk(clk),
	.d(\addr_cmd~519_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr0),
	.prn(vcc));
defparam \addr_cmd[0].addr[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[0] .power_up = "low";

dffeas \addr_cmd[0].addr[1] (
	.clk(clk),
	.d(\addr_cmd~523_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr1),
	.prn(vcc));
defparam \addr_cmd[0].addr[1] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[1] .power_up = "low";

dffeas \addr_cmd[0].addr[4] (
	.clk(clk),
	.d(\addr_cmd~524_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr4),
	.prn(vcc));
defparam \addr_cmd[0].addr[4] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[4] .power_up = "low";

dffeas \addr_cmd[0].addr[8] (
	.clk(clk),
	.d(\addr_cmd~526_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr8),
	.prn(vcc));
defparam \addr_cmd[0].addr[8] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[8] .power_up = "low";

dffeas \addr_cmd[0].addr[10] (
	.clk(clk),
	.d(\addr_cmd~531_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr10),
	.prn(vcc));
defparam \addr_cmd[0].addr[10] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[10] .power_up = "low";

dffeas \addr_cmd[0].ba[0] (
	.clk(clk),
	.d(\addr_cmd~535_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ba0),
	.prn(vcc));
defparam \addr_cmd[0].ba[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].ba[0] .power_up = "low";

dffeas \addr_cmd[0].ba[1] (
	.clk(clk),
	.d(\addr_cmd~537_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ba1),
	.prn(vcc));
defparam \addr_cmd[0].ba[1] .is_wysiwyg = "true";
defparam \addr_cmd[0].ba[1] .power_up = "low";

dffeas \addr_cmd[0].ras_n (
	.clk(clk),
	.d(\addr_cmd~538_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ras_n),
	.prn(vcc));
defparam \addr_cmd[0].ras_n .is_wysiwyg = "true";
defparam \addr_cmd[0].ras_n .power_up = "low";

dffeas \addr_cmd[0].cas_n (
	.clk(clk),
	.d(\addr_cmd~549_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0cas_n),
	.prn(vcc));
defparam \addr_cmd[0].cas_n .is_wysiwyg = "true";
defparam \addr_cmd[0].cas_n .power_up = "low";

dffeas \addr_cmd[0].we_n (
	.clk(clk),
	.d(\addr_cmd~550_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0we_n),
	.prn(vcc));
defparam \addr_cmd[0].we_n .is_wysiwyg = "true";
defparam \addr_cmd[0].we_n .power_up = "low";

dffeas \admin_ctrl.command_done (
	.clk(clk),
	.d(\command_done~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(admin_ctrlcommand_done),
	.prn(vcc));
defparam \admin_ctrl.command_done .is_wysiwyg = "true";
defparam \admin_ctrl.command_done .power_up = "low";

cycloneiii_lcell_comb \state~172 (
	.dataa(\state.s_access~q ),
	.datab(dgwb_ac_access_req),
	.datac(dgrb_ac_access_req),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~172_combout ),
	.cout());
defparam \state~172 .lut_mask = 16'hBEBE;
defparam \state~172 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~168 (
	.dataa(\state.s_idle~q ),
	.datab(dgwb_ac_access_req),
	.datac(dgrb_ac_access_req),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~168_combout ),
	.cout());
defparam \state~168 .lut_mask = 16'hBEBE;
defparam \state~168 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector15~0 (
	.dataa(\Selector10~1_combout ),
	.datab(\process_10~0_combout ),
	.datac(\state~168_combout ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hFEFF;
defparam \Selector15~0 .sum_lutc_input = "datac";

dffeas command_started(
	.clk(clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\command_started~q ),
	.prn(vcc));
defparam command_started.is_wysiwyg = "true";
defparam command_started.power_up = "low";

cycloneiii_lcell_comb \admin_req_extended~2 (
	.dataa(ac_muxctrl_broadcast_rcommand_req),
	.datab(\admin_req_extended~q ),
	.datac(Selector1),
	.datad(\command_started~q ),
	.cin(gnd),
	.combout(\admin_req_extended~2_combout ),
	.cout());
defparam \admin_req_extended~2 .lut_mask = 16'hEFFF;
defparam \admin_req_extended~2 .sum_lutc_input = "datac";

dffeas admin_req_extended(
	.clk(clk),
	.d(\admin_req_extended~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\admin_req_extended~q ),
	.prn(vcc));
defparam admin_req_extended.is_wysiwyg = "true";
defparam admin_req_extended.power_up = "low";

cycloneiii_lcell_comb \process_10~0 (
	.dataa(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datab(\admin_req_extended~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_10~0_combout ),
	.cout());
defparam \process_10~0 .lut_mask = 16'hEEEE;
defparam \process_10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~173 (
	.dataa(\state~171_combout ),
	.datab(\state~172_combout ),
	.datac(\process_10~0_combout ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\state~173_combout ),
	.cout());
defparam \state~173 .lut_mask = 16'hFEFF;
defparam \state~173 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~175 (
	.dataa(ctl_init_success),
	.datab(gnd),
	.datac(\state.s_reset~q ),
	.datad(\state~173_combout ),
	.cin(gnd),
	.combout(\state~175_combout ),
	.cout());
defparam \state~175 .lut_mask = 16'hFFF5;
defparam \state~175 .sum_lutc_input = "datac";

dffeas \state.s_reset (
	.clk(clk),
	.d(\state~175_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_reset~q ),
	.prn(vcc));
defparam \state.s_reset .is_wysiwyg = "true";
defparam \state.s_reset .power_up = "low";

cycloneiii_lcell_comb \state~177 (
	.dataa(\state~176_combout ),
	.datab(\state.s_run_init_seq~q ),
	.datac(\state~173_combout ),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\state~177_combout ),
	.cout());
defparam \state~177 .lut_mask = 16'hACFF;
defparam \state~177 .sum_lutc_input = "datac";

dffeas \state.s_run_init_seq (
	.clk(clk),
	.d(\state~177_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_run_init_seq~q ),
	.prn(vcc));
defparam \state.s_run_init_seq .is_wysiwyg = "true";
defparam \state.s_run_init_seq .power_up = "low";

cycloneiii_lcell_comb \addr_cmd[0].cke[0]~0 (
	.dataa(\state.s_reset~q ),
	.datab(addr_cmd0cke0),
	.datac(gnd),
	.datad(\state.s_run_init_seq~q ),
	.cin(gnd),
	.combout(\addr_cmd[0].cke[0]~0_combout ),
	.cout());
defparam \addr_cmd[0].cke[0]~0 .lut_mask = 16'hAACC;
defparam \addr_cmd[0].cke[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector286~2 (
	.dataa(\ac_state.s_10~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.s_run_init_seq~q ),
	.cin(gnd),
	.combout(\Selector286~2_combout ),
	.cout());
defparam \Selector286~2 .lut_mask = 16'hAAFF;
defparam \Selector286~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector2~1 (
	.dataa(\Selector2~0_combout ),
	.datab(\state.s_run_init_seq~q ),
	.datac(\finished_state~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFEFE;
defparam \Selector2~1 .sum_lutc_input = "datac";

dffeas \state.s_program_cal_mrs (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_program_cal_mrs~q ),
	.prn(vcc));
defparam \state.s_program_cal_mrs .is_wysiwyg = "true";
defparam \state.s_program_cal_mrs .power_up = "low";

cycloneiii_lcell_comb \WideOr41~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_run_init_seq~q ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\WideOr41~0_combout ),
	.cout());
defparam \WideOr41~0 .lut_mask = 16'h0FFF;
defparam \WideOr41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_7~0 (
	.dataa(\Equal0~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\process_7~0_combout ),
	.cout());
defparam \process_7~0 .lut_mask = 16'hAAFF;
defparam \process_7~0 .sum_lutc_input = "datac";

dffeas refresh_due(
	.clk(clk),
	.d(\process_7~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_due~q ),
	.prn(vcc));
defparam refresh_due.is_wysiwyg = "true";
defparam refresh_due.power_up = "low";

cycloneiii_lcell_comb \process_8~4 (
	.dataa(\num_stacked_refreshes[2]~q ),
	.datab(\num_stacked_refreshes[1]~q ),
	.datac(\num_stacked_refreshes[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_8~4_combout ),
	.cout());
defparam \process_8~4 .lut_mask = 16'hFEFE;
defparam \process_8~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \num_stacked_refreshes~13 (
	.dataa(\refresh_due~q ),
	.datab(\process_8~4_combout ),
	.datac(\process_8~1_combout ),
	.datad(\num_stacked_refreshes[0]~q ),
	.cin(gnd),
	.combout(\num_stacked_refreshes~13_combout ),
	.cout());
defparam \num_stacked_refreshes~13 .lut_mask = 16'h6996;
defparam \num_stacked_refreshes~13 .sum_lutc_input = "datac";

dffeas \num_stacked_refreshes[0] (
	.clk(clk),
	.d(\num_stacked_refreshes~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[0]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[0] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[0] .power_up = "low";

cycloneiii_lcell_comb \process_8~1 (
	.dataa(\refresh_done~q ),
	.datab(\num_stacked_refreshes[2]~q ),
	.datac(\num_stacked_refreshes[1]~q ),
	.datad(\num_stacked_refreshes[0]~q ),
	.cin(gnd),
	.combout(\process_8~1_combout ),
	.cout());
defparam \process_8~1 .lut_mask = 16'hBFFF;
defparam \process_8~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \num_stacked_refreshes~11 (
	.dataa(\num_stacked_refreshes[0]~q ),
	.datab(\refresh_due~q ),
	.datac(\process_8~1_combout ),
	.datad(\process_8~4_combout ),
	.cin(gnd),
	.combout(\num_stacked_refreshes~11_combout ),
	.cout());
defparam \num_stacked_refreshes~11 .lut_mask = 16'h6FFF;
defparam \num_stacked_refreshes~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \num_stacked_refreshes~12 (
	.dataa(ctl_init_success),
	.datab(gnd),
	.datac(\num_stacked_refreshes[1]~q ),
	.datad(\num_stacked_refreshes~11_combout ),
	.cin(gnd),
	.combout(\num_stacked_refreshes~12_combout ),
	.cout());
defparam \num_stacked_refreshes~12 .lut_mask = 16'h5FF5;
defparam \num_stacked_refreshes~12 .sum_lutc_input = "datac";

dffeas \num_stacked_refreshes[1] (
	.clk(clk),
	.d(\num_stacked_refreshes~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[1]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[1] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[1] .power_up = "low";

cycloneiii_lcell_comb \Selector3~3 (
	.dataa(\state.s_refresh_done~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'hEEEE;
defparam \Selector3~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~1 (
	.dataa(dgwb_ac_access_req),
	.datab(dgrb_ac_access_req),
	.datac(curr_cmdcmd_prep_customer_mr_setup),
	.datad(\admin_req_extended~q ),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'h6FFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~4 (
	.dataa(\refreshes_maxed~q ),
	.datab(\Selector3~3_combout ),
	.datac(\state.s_topup_refresh_done~q ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
defparam \Selector3~4 .lut_mask = 16'hFFFE;
defparam \Selector3~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~178 (
	.dataa(\state~172_combout ),
	.datab(\state.s_access_precharge~q ),
	.datac(\state~173_combout ),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\state~178_combout ),
	.cout());
defparam \state~178 .lut_mask = 16'hACFF;
defparam \state~178 .sum_lutc_input = "datac";

dffeas \state.s_access_precharge (
	.clk(clk),
	.d(\state~178_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access_precharge~q ),
	.prn(vcc));
defparam \state.s_access_precharge .is_wysiwyg = "true";
defparam \state.s_access_precharge .power_up = "low";

cycloneiii_lcell_comb \Selector3~5 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\state.s_access_precharge~q ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(\mem_init_complete~q ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
defparam \Selector3~5 .lut_mask = 16'hFEFF;
defparam \Selector3~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector3~6 (
	.dataa(\Selector3~2_combout ),
	.datab(\finished_state~q ),
	.datac(\Selector3~4_combout ),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
defparam \Selector3~6 .lut_mask = 16'hFFFE;
defparam \Selector3~6 .sum_lutc_input = "datac";

dffeas \state.s_idle (
	.clk(clk),
	.d(\Selector3~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_idle~q ),
	.prn(vcc));
defparam \state.s_idle .is_wysiwyg = "true";
defparam \state.s_idle .power_up = "low";

cycloneiii_lcell_comb \Selector216~0 (
	.dataa(\state.s_access~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\state.s_idle~q ),
	.datad(\state.s_run_init_seq~q ),
	.cin(gnd),
	.combout(\Selector216~0_combout ),
	.cout());
defparam \Selector216~0 .lut_mask = 16'hFEFF;
defparam \Selector216~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector216~1 (
	.dataa(\ac_state.s_8~q ),
	.datab(\per_cs_init_seen[0]~q ),
	.datac(\Selector216~0_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\Selector216~1_combout ),
	.cout());
defparam \Selector216~1 .lut_mask = 16'hFFFE;
defparam \Selector216~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~28 (
	.dataa(\stage_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~27 ),
	.combout(\Add3~28_combout ),
	.cout(\Add3~29 ));
defparam \Add3~28 .lut_mask = 16'h5A5F;
defparam \Add3~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~30 (
	.dataa(\stage_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~29 ),
	.combout(\Add3~30_combout ),
	.cout(\Add3~31 ));
defparam \Add3~30 .lut_mask = 16'h5AAF;
defparam \Add3~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~32 (
	.dataa(\stage_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~31 ),
	.combout(\Add3~32_combout ),
	.cout(\Add3~33 ));
defparam \Add3~32 .lut_mask = 16'h5A5F;
defparam \Add3~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~38 (
	.dataa(\stage_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~37 ),
	.combout(\Add3~38_combout ),
	.cout(\Add3~39 ));
defparam \Add3~38 .lut_mask = 16'h5AAF;
defparam \Add3~38 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~40 (
	.dataa(\stage_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~39 ),
	.combout(\Add3~40_combout ),
	.cout(\Add3~41 ));
defparam \Add3~40 .lut_mask = 16'h5A5F;
defparam \Add3~40 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add3~94 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~94_combout ),
	.cout());
defparam \Add3~94 .lut_mask = 16'hFEFE;
defparam \Add3~94 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~1 (
	.dataa(gnd),
	.datab(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datac(\admin_req_extended~q ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
defparam \Selector8~1 .lut_mask = 16'h3FFF;
defparam \Selector8~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector8~2 (
	.dataa(\Selector8~0_combout ),
	.datab(\state.s_access~q ),
	.datac(dgb_ac_access_req),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
defparam \Selector8~2 .lut_mask = 16'hFFFE;
defparam \Selector8~2 .sum_lutc_input = "datac";

dffeas \state.s_access (
	.clk(clk),
	.d(\Selector8~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access~q ),
	.prn(vcc));
defparam \state.s_access .is_wysiwyg = "true";
defparam \state.s_access .power_up = "low";

cycloneiii_lcell_comb \state~166 (
	.dataa(\state.s_reset~q ),
	.datab(gnd),
	.datac(\state.s_access~q ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\state~166_combout ),
	.cout());
defparam \state~166 .lut_mask = 16'hAFFF;
defparam \state~166 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state.s_10~5 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\state~166_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\ac_state.s_10~5_combout ),
	.cout());
defparam \ac_state.s_10~5 .lut_mask = 16'hF7FF;
defparam \ac_state.s_10~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state.s_10~3 (
	.dataa(\process_12~6_combout ),
	.datab(\ac_state.s_10~5_combout ),
	.datac(\state~166_combout ),
	.datad(\WideOr41~0_combout ),
	.cin(gnd),
	.combout(\ac_state.s_10~3_combout ),
	.cout());
defparam \ac_state.s_10~3 .lut_mask = 16'hEFFF;
defparam \ac_state.s_10~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state.s_10~4 (
	.dataa(\ac_state.s_9~q ),
	.datab(\ac_state.s_10~3_combout ),
	.datac(\ac_state.s_10~q ),
	.datad(\ac_state.s_10~5_combout ),
	.cin(gnd),
	.combout(\ac_state.s_10~4_combout ),
	.cout());
defparam \ac_state.s_10~4 .lut_mask = 16'hFEFF;
defparam \ac_state.s_10~4 .sum_lutc_input = "datac";

dffeas \ac_state.s_10 (
	.clk(clk),
	.d(\ac_state.s_10~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_10~q ),
	.prn(vcc));
defparam \ac_state.s_10 .is_wysiwyg = "true";
defparam \ac_state.s_10 .power_up = "low";

cycloneiii_lcell_comb \Selector228~1 (
	.dataa(\Selector228~0_combout ),
	.datab(\ac_state.s_11~q ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(\state~166_combout ),
	.cin(gnd),
	.combout(\Selector228~1_combout ),
	.cout());
defparam \Selector228~1 .lut_mask = 16'hFEFF;
defparam \Selector228~1 .sum_lutc_input = "datac";

dffeas \ac_state.s_11 (
	.clk(clk),
	.d(\Selector228~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_12~2_combout ),
	.q(\ac_state.s_11~q ),
	.prn(vcc));
defparam \ac_state.s_11 .is_wysiwyg = "true";
defparam \ac_state.s_11 .power_up = "low";

cycloneiii_lcell_comb \WideOr38~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_access~q ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\WideOr38~1_combout ),
	.cout());
defparam \WideOr38~1 .lut_mask = 16'h0FFF;
defparam \WideOr38~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr41~1 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\state.s_reset~q ),
	.datad(\WideOr38~1_combout ),
	.cin(gnd),
	.combout(\WideOr41~1_combout ),
	.cout());
defparam \WideOr41~1 .lut_mask = 16'hEFFF;
defparam \WideOr41~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~90 (
	.dataa(\ac_state.s_8~q ),
	.datab(\WideOr41~1_combout ),
	.datac(\process_12~6_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\ac_state~90_combout ),
	.cout());
defparam \ac_state~90 .lut_mask = 16'hFFFE;
defparam \ac_state~90 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~91 (
	.dataa(\state.s_access~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\state.s_idle~q ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\ac_state~91_combout ),
	.cout());
defparam \ac_state~91 .lut_mask = 16'hFF7F;
defparam \ac_state~91 .sum_lutc_input = "datac";

dffeas \ac_state.s_9 (
	.clk(clk),
	.d(\ac_state~90_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_9~q ),
	.prn(vcc));
defparam \ac_state.s_9 .is_wysiwyg = "true";
defparam \ac_state.s_9 .power_up = "low";

cycloneiii_lcell_comb \WideOr26~0 (
	.dataa(gnd),
	.datab(\ac_state.s_10~q ),
	.datac(\ac_state.s_9~q ),
	.datad(\ac_state.s_11~q ),
	.cin(gnd),
	.combout(\WideOr26~0_combout ),
	.cout());
defparam \WideOr26~0 .lut_mask = 16'h3FFF;
defparam \WideOr26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \finished_state~1 (
	.dataa(\ac_state.s_9~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\finished_state~1_combout ),
	.cout());
defparam \finished_state~1 .lut_mask = 16'hEEEE;
defparam \finished_state~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector217~2 (
	.dataa(\Selector217~1_combout ),
	.datab(\finished_state~1_combout ),
	.datac(\ac_state.s_0~q ),
	.datad(\state~166_combout ),
	.cin(gnd),
	.combout(\Selector217~2_combout ),
	.cout());
defparam \Selector217~2 .lut_mask = 16'hEFFF;
defparam \Selector217~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector286~3 (
	.dataa(\ac_state.s_11~q ),
	.datab(gnd),
	.datac(\ac_state.s_10~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\Selector286~3_combout ),
	.cout());
defparam \Selector286~3 .lut_mask = 16'hAFFF;
defparam \Selector286~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector217~3 (
	.dataa(\Selector217~0_combout ),
	.datab(\Selector217~2_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\Selector286~3_combout ),
	.cin(gnd),
	.combout(\Selector217~3_combout ),
	.cout());
defparam \Selector217~3 .lut_mask = 16'h7FFF;
defparam \Selector217~3 .sum_lutc_input = "datac";

dffeas \ac_state.s_0 (
	.clk(clk),
	.d(\Selector217~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_12~2_combout ),
	.q(\ac_state.s_0~q ),
	.prn(vcc));
defparam \ac_state.s_0 .is_wysiwyg = "true";
defparam \ac_state.s_0 .power_up = "low";

cycloneiii_lcell_comb \process_10~1 (
	.dataa(curr_cmdcmd_prep_customer_mr_setup),
	.datab(\admin_req_extended~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_10~1_combout ),
	.cout());
defparam \process_10~1 .lut_mask = 16'hEEEE;
defparam \process_10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~1 (
	.dataa(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datab(\admin_req_extended~q ),
	.datac(\state.s_reset~q ),
	.datad(\finished_state~q ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'h7FFF;
defparam \Selector7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector10~0 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\process_10~1_combout ),
	.datac(\Selector7~0_combout ),
	.datad(\Selector7~1_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFFFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

dffeas \state.s_prog_user_mrs (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_prog_user_mrs~q ),
	.prn(vcc));
defparam \state.s_prog_user_mrs .is_wysiwyg = "true";
defparam \state.s_prog_user_mrs .power_up = "low";

cycloneiii_lcell_comb \ac_state~93 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\state~166_combout ),
	.datad(\state.s_run_init_seq~q ),
	.cin(gnd),
	.combout(\ac_state~93_combout ),
	.cout());
defparam \ac_state~93 .lut_mask = 16'hEFFF;
defparam \ac_state~93 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~94 (
	.dataa(\ac_state.s_6~q ),
	.datab(\ac_state~93_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\ac_state~94_combout ),
	.cout());
defparam \ac_state~94 .lut_mask = 16'hFFFE;
defparam \ac_state~94 .sum_lutc_input = "datac";

dffeas \ac_state.s_7 (
	.clk(clk),
	.d(\ac_state~94_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_7~q ),
	.prn(vcc));
defparam \ac_state.s_7 .is_wysiwyg = "true";
defparam \ac_state.s_7 .power_up = "low";

cycloneiii_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_2~q ),
	.datad(\ac_state.s_7~q ),
	.cin(gnd),
	.combout(\Add3~21_combout ),
	.cout());
defparam \Add3~21 .lut_mask = 16'h0FFF;
defparam \Add3~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~95 (
	.dataa(\ac_state.s_5~q ),
	.datab(\ac_state~93_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\ac_state~95_combout ),
	.cout());
defparam \ac_state~95 .lut_mask = 16'hFFFE;
defparam \ac_state~95 .sum_lutc_input = "datac";

dffeas \ac_state.s_6 (
	.clk(clk),
	.d(\ac_state~95_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_6~q ),
	.prn(vcc));
defparam \ac_state.s_6 .is_wysiwyg = "true";
defparam \ac_state.s_6 .power_up = "low";

cycloneiii_lcell_comb \ac_state~97 (
	.dataa(\ac_state.s_4~q ),
	.datab(\ac_state~93_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\ac_state~97_combout ),
	.cout());
defparam \ac_state~97 .lut_mask = 16'hFFFE;
defparam \ac_state~97 .sum_lutc_input = "datac";

dffeas \ac_state.s_5 (
	.clk(clk),
	.d(\ac_state~97_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_5~q ),
	.prn(vcc));
defparam \ac_state.s_5 .is_wysiwyg = "true";
defparam \ac_state.s_5 .power_up = "low";

cycloneiii_lcell_comb \process_12~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_6~q ),
	.datad(\ac_state.s_5~q ),
	.cin(gnd),
	.combout(\process_12~4_combout ),
	.cout());
defparam \process_12~4 .lut_mask = 16'h0FFF;
defparam \process_12~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~92 (
	.dataa(\ac_state.s_7~q ),
	.datab(\WideOr41~1_combout ),
	.datac(\process_12~6_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\ac_state~92_combout ),
	.cout());
defparam \ac_state~92 .lut_mask = 16'hFFFE;
defparam \ac_state~92 .sum_lutc_input = "datac";

dffeas \ac_state.s_8 (
	.clk(clk),
	.d(\ac_state~92_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_8~q ),
	.prn(vcc));
defparam \ac_state.s_8 .is_wysiwyg = "true";
defparam \ac_state.s_8 .power_up = "low";

cycloneiii_lcell_comb \process_12~5 (
	.dataa(\Add3~20_combout ),
	.datab(\Add3~21_combout ),
	.datac(\process_12~4_combout ),
	.datad(\ac_state.s_8~q ),
	.cin(gnd),
	.combout(\process_12~5_combout ),
	.cout());
defparam \process_12~5 .lut_mask = 16'hFEFF;
defparam \process_12~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_12~6 (
	.dataa(\ac_state.s_9~q ),
	.datab(\WideOr26~0_combout ),
	.datac(\ac_state.s_0~q ),
	.datad(\process_12~5_combout ),
	.cin(gnd),
	.combout(\process_12~6_combout ),
	.cout());
defparam \process_12~6 .lut_mask = 16'hEFFE;
defparam \process_12~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~121 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\ac_state.s_10~q ),
	.datac(\ac_state.s_11~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\stage_counter[17]~121_combout ),
	.cout());
defparam \stage_counter[17]~121 .lut_mask = 16'hBFFF;
defparam \stage_counter[17]~121 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~118 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\stage_counter[17]~118_combout ),
	.cout());
defparam \stage_counter[17]~118 .lut_mask = 16'hFFF0;
defparam \stage_counter[17]~118 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~6 (
	.dataa(gnd),
	.datab(\state.s_topup_refresh~q ),
	.datac(\state.s_refresh~q ),
	.datad(\state.s_access_act~q ),
	.cin(gnd),
	.combout(\Selector269~6_combout ),
	.cout());
defparam \Selector269~6 .lut_mask = 16'h3FFF;
defparam \Selector269~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~123 (
	.dataa(\WideNor1~0_combout ),
	.datab(\state.s_access_precharge~q ),
	.datac(\Selector269~6_combout ),
	.datad(\ac_state.s_2~q ),
	.cin(gnd),
	.combout(\stage_counter[17]~123_combout ),
	.cout());
defparam \stage_counter[17]~123 .lut_mask = 16'hEFFF;
defparam \stage_counter[17]~123 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state.s_1~1 (
	.dataa(\ac_state.s_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac_state.s_1~1_combout ),
	.cout());
defparam \ac_state.s_1~1 .lut_mask = 16'h5555;
defparam \ac_state.s_1~1 .sum_lutc_input = "datac";

dffeas \ac_state.s_1 (
	.clk(clk),
	.d(\ac_state.s_1~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_1~q ),
	.prn(vcc));
defparam \ac_state.s_1 .is_wysiwyg = "true";
defparam \ac_state.s_1 .power_up = "low";

cycloneiii_lcell_comb \state~174 (
	.dataa(\state~169_combout ),
	.datab(\state.s_dummy_wait~q ),
	.datac(\state~173_combout ),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\state~174_combout ),
	.cout());
defparam \state~174 .lut_mask = 16'hACFF;
defparam \state~174 .sum_lutc_input = "datac";

dffeas \state.s_dummy_wait (
	.clk(clk),
	.d(\state~174_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_dummy_wait~q ),
	.prn(vcc));
defparam \state.s_dummy_wait .is_wysiwyg = "true";
defparam \state.s_dummy_wait .power_up = "low";

cycloneiii_lcell_comb \WideOr45~1 (
	.dataa(gnd),
	.datab(\state.s_dummy_wait~q ),
	.datac(\state.s_topup_refresh_done~q ),
	.datad(\state.s_refresh_done~q ),
	.cin(gnd),
	.combout(\WideOr45~1_combout ),
	.cout());
defparam \WideOr45~1 .lut_mask = 16'h3FFF;
defparam \WideOr45~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~139 (
	.dataa(\ac_state.s_0~q ),
	.datab(\ac_state.s_1~q ),
	.datac(\WideOr45~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter[17]~139_combout ),
	.cout());
defparam \stage_counter[17]~139 .lut_mask = 16'hBFBF;
defparam \stage_counter[17]~139 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~124 (
	.dataa(\stage_counter[17]~122_combout ),
	.datab(\stage_counter[17]~118_combout ),
	.datac(\stage_counter[17]~123_combout ),
	.datad(\stage_counter[17]~139_combout ),
	.cin(gnd),
	.combout(\stage_counter[17]~124_combout ),
	.cout());
defparam \stage_counter[17]~124 .lut_mask = 16'hFFFB;
defparam \stage_counter[17]~124 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[17]~125 (
	.dataa(\stage_counter[17]~120_combout ),
	.datab(\stage_counter[17]~121_combout ),
	.datac(\stage_counter[17]~124_combout ),
	.datad(\state.s_run_init_seq~q ),
	.cin(gnd),
	.combout(\stage_counter[17]~125_combout ),
	.cout());
defparam \stage_counter[17]~125 .lut_mask = 16'hFF7F;
defparam \stage_counter[17]~125 .sum_lutc_input = "datac";

dffeas \stage_counter[10] (
	.clk(clk),
	.d(\Add3~94_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[10]~q ),
	.prn(vcc));
defparam \stage_counter[10] .is_wysiwyg = "true";
defparam \stage_counter[10] .power_up = "low";

cycloneiii_lcell_comb \Add3~95 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~95_combout ),
	.cout());
defparam \Add3~95 .lut_mask = 16'hFEFE;
defparam \Add3~95 .sum_lutc_input = "datac";

dffeas \stage_counter[9] (
	.clk(clk),
	.d(\Add3~95_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[9]~q ),
	.prn(vcc));
defparam \stage_counter[9] .is_wysiwyg = "true";
defparam \stage_counter[9] .power_up = "low";

cycloneiii_lcell_comb \Add3~96 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter_zero~q ),
	.datac(\Add3~38_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~96_combout ),
	.cout());
defparam \Add3~96 .lut_mask = 16'hFEFE;
defparam \Add3~96 .sum_lutc_input = "datac";

dffeas \stage_counter[8] (
	.clk(clk),
	.d(\Add3~96_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~125_combout ),
	.q(\stage_counter[8]~q ),
	.prn(vcc));
defparam \stage_counter[8] .is_wysiwyg = "true";
defparam \stage_counter[8] .power_up = "low";

cycloneiii_lcell_comb \stage_counter_zero~3 (
	.dataa(\stage_counter[11]~q ),
	.datab(\stage_counter[10]~q ),
	.datac(\stage_counter[9]~q ),
	.datad(\stage_counter[8]~q ),
	.cin(gnd),
	.combout(\stage_counter_zero~3_combout ),
	.cout());
defparam \stage_counter_zero~3 .lut_mask = 16'h7FFF;
defparam \stage_counter_zero~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb WideOr26(
	.dataa(\ac_state.s_10~q ),
	.datab(\ac_state.s_9~q ),
	.datac(\ac_state.s_8~q ),
	.datad(\ac_state.s_11~q ),
	.cin(gnd),
	.combout(\WideOr26~combout ),
	.cout());
defparam WideOr26.lut_mask = 16'hFFFE;
defparam WideOr26.sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~126 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\WideOr26~combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter[5]~126_combout ),
	.cout());
defparam \stage_counter[5]~126 .lut_mask = 16'hEEEE;
defparam \stage_counter[5]~126 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~61 (
	.dataa(\WideOr26~1_combout ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\stage_counter[17]~123_combout ),
	.datad(\stage_counter[5]~126_combout ),
	.cin(gnd),
	.combout(\Add3~61_combout ),
	.cout());
defparam \Add3~61 .lut_mask = 16'hBFFF;
defparam \Add3~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~62 (
	.dataa(\Add3~60_combout ),
	.datab(\stage_counter[17]~121_combout ),
	.datac(\stage_counter[17]~139_combout ),
	.datad(\Add3~61_combout ),
	.cin(gnd),
	.combout(\Add3~62_combout ),
	.cout());
defparam \Add3~62 .lut_mask = 16'hFEFF;
defparam \Add3~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~65 (
	.dataa(\Add3~64_combout ),
	.datab(\stage_counter[6]~q ),
	.datac(\Add3~62_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~65_combout ),
	.cout());
defparam \Add3~65 .lut_mask = 16'hFEFE;
defparam \Add3~65 .sum_lutc_input = "datac";

dffeas \stage_counter[6] (
	.clk(clk),
	.d(\Add3~65_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[6]~q ),
	.prn(vcc));
defparam \stage_counter[6] .is_wysiwyg = "true";
defparam \stage_counter[6] .power_up = "low";

cycloneiii_lcell_comb \stage_counter~127 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter~127_combout ),
	.cout());
defparam \stage_counter~127 .lut_mask = 16'hEEEE;
defparam \stage_counter~127 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector19~0 (
	.dataa(\ac_state.s_10~q ),
	.datab(\stage_counter~127_combout ),
	.datac(\ac_state.s_11~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
defparam \Selector19~0 .lut_mask = 16'hEFFF;
defparam \Selector19~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~129 (
	.dataa(\ac_state.s_0~q ),
	.datab(\state.s_dummy_wait~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\state.s_prog_user_mrs~q ),
	.cin(gnd),
	.combout(\stage_counter[5]~129_combout ),
	.cout());
defparam \stage_counter[5]~129 .lut_mask = 16'hEFFF;
defparam \stage_counter[5]~129 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~130 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_refresh_done~q ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\stage_counter[5]~130_combout ),
	.cout());
defparam \stage_counter[5]~130 .lut_mask = 16'hFEFF;
defparam \stage_counter[5]~130 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~131 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_refresh_done~q ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter[5]~131_combout ),
	.cout());
defparam \stage_counter[5]~131 .lut_mask = 16'hFEFE;
defparam \stage_counter[5]~131 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter[5]~132 (
	.dataa(\stage_counter[5]~128_combout ),
	.datab(\stage_counter[5]~129_combout ),
	.datac(\stage_counter[5]~130_combout ),
	.datad(\stage_counter[5]~131_combout ),
	.cin(gnd),
	.combout(\stage_counter[5]~132_combout ),
	.cout());
defparam \stage_counter[5]~132 .lut_mask = 16'hFEFF;
defparam \stage_counter[5]~132 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector192~0 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[5]~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Selector192~0_combout ),
	.cout());
defparam \Selector192~0 .lut_mask = 16'hEFFF;
defparam \Selector192~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter~133 (
	.dataa(\Selector37~0_combout ),
	.datab(\Selector192~0_combout ),
	.datac(\stage_counter[5]~131_combout ),
	.datad(\stage_counter[5]~130_combout ),
	.cin(gnd),
	.combout(\stage_counter~133_combout ),
	.cout());
defparam \stage_counter~133 .lut_mask = 16'hEFFE;
defparam \stage_counter~133 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter~134 (
	.dataa(\stage_counter~127_combout ),
	.datab(\Selector19~0_combout ),
	.datac(\stage_counter[5]~132_combout ),
	.datad(\stage_counter~133_combout ),
	.cin(gnd),
	.combout(\stage_counter~134_combout ),
	.cout());
defparam \stage_counter~134 .lut_mask = 16'hEFFE;
defparam \stage_counter~134 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~66 (
	.dataa(\state~166_combout ),
	.datab(\stage_counter~134_combout ),
	.datac(\Add3~32_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~66_combout ),
	.cout());
defparam \Add3~66 .lut_mask = 16'hFAFC;
defparam \Add3~66 .sum_lutc_input = "datac";

dffeas \stage_counter[5] (
	.clk(clk),
	.d(\Add3~66_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[5]~q ),
	.prn(vcc));
defparam \stage_counter[5] .is_wysiwyg = "true";
defparam \stage_counter[5] .power_up = "low";

cycloneiii_lcell_comb \stage_counter~135 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stage_counter~135_combout ),
	.cout());
defparam \stage_counter~135 .lut_mask = 16'hEEEE;
defparam \stage_counter~135 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector20~0 (
	.dataa(\process_12~6_combout ),
	.datab(\stage_counter~135_combout ),
	.datac(\ac_state.s_10~q ),
	.datad(\ac_state.s_11~q ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'hEFFF;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector193~0 (
	.dataa(\state.s_reset~q ),
	.datab(\stage_counter[4]~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Selector193~0_combout ),
	.cout());
defparam \Selector193~0 .lut_mask = 16'hEFFF;
defparam \Selector193~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter~136 (
	.dataa(\Selector38~0_combout ),
	.datab(\Selector193~0_combout ),
	.datac(\stage_counter[5]~131_combout ),
	.datad(\stage_counter[5]~130_combout ),
	.cin(gnd),
	.combout(\stage_counter~136_combout ),
	.cout());
defparam \stage_counter~136 .lut_mask = 16'hEFFE;
defparam \stage_counter~136 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter~137 (
	.dataa(\stage_counter~135_combout ),
	.datab(\Selector20~0_combout ),
	.datac(\stage_counter[5]~132_combout ),
	.datad(\stage_counter~136_combout ),
	.cin(gnd),
	.combout(\stage_counter~137_combout ),
	.cout());
defparam \stage_counter~137 .lut_mask = 16'hEFFE;
defparam \stage_counter~137 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~67 (
	.dataa(\state~166_combout ),
	.datab(\stage_counter~137_combout ),
	.datac(\Add3~30_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~67_combout ),
	.cout());
defparam \Add3~67 .lut_mask = 16'hFAFC;
defparam \Add3~67 .sum_lutc_input = "datac";

dffeas \stage_counter[4] (
	.clk(clk),
	.d(\Add3~67_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[4]~q ),
	.prn(vcc));
defparam \stage_counter[4] .is_wysiwyg = "true";
defparam \stage_counter[4] .power_up = "low";

cycloneiii_lcell_comb \stage_counter_zero~4 (
	.dataa(\stage_counter[7]~q ),
	.datab(\stage_counter[6]~q ),
	.datac(\stage_counter[5]~q ),
	.datad(\stage_counter[4]~q ),
	.cin(gnd),
	.combout(\stage_counter_zero~4_combout ),
	.cout());
defparam \stage_counter_zero~4 .lut_mask = 16'h7FFF;
defparam \stage_counter_zero~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~70 (
	.dataa(\state.s_access_precharge~q ),
	.datab(\state.s_reset~q ),
	.datac(\stage_counter_zero~q ),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Add3~70_combout ),
	.cout());
defparam \Add3~70 .lut_mask = 16'hBFFF;
defparam \Add3~70 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~71 (
	.dataa(\addr_cmd~521_combout ),
	.datab(\Add3~70_combout ),
	.datac(\Add3~28_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\Add3~71_combout ),
	.cout());
defparam \Add3~71 .lut_mask = 16'hFEFF;
defparam \Add3~71 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~72 (
	.dataa(\Add3~69_combout ),
	.datab(\Add3~71_combout ),
	.datac(\stage_counter[3]~q ),
	.datad(\Add3~62_combout ),
	.cin(gnd),
	.combout(\Add3~72_combout ),
	.cout());
defparam \Add3~72 .lut_mask = 16'hFFFE;
defparam \Add3~72 .sum_lutc_input = "datac";

dffeas \stage_counter[3] (
	.clk(clk),
	.d(\Add3~72_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[3]~q ),
	.prn(vcc));
defparam \stage_counter[3] .is_wysiwyg = "true";
defparam \stage_counter[3] .power_up = "low";

cycloneiii_lcell_comb \Add3~60 (
	.dataa(\state.s_reset~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\Add3~60_combout ),
	.cout());
defparam \Add3~60 .lut_mask = 16'hAAFF;
defparam \Add3~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~79 (
	.dataa(\stage_counter[17]~121_combout ),
	.datab(\ac_state.s_1~q ),
	.datac(\WideOr45~1_combout ),
	.datad(\Add3~61_combout ),
	.cin(gnd),
	.combout(\Add3~79_combout ),
	.cout());
defparam \Add3~79 .lut_mask = 16'hBFFF;
defparam \Add3~79 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~80 (
	.dataa(\Add3~78_combout ),
	.datab(\stage_counter[2]~q ),
	.datac(\Add3~60_combout ),
	.datad(\Add3~79_combout ),
	.cin(gnd),
	.combout(\Add3~80_combout ),
	.cout());
defparam \Add3~80 .lut_mask = 16'hFFFE;
defparam \Add3~80 .sum_lutc_input = "datac";

dffeas \stage_counter[2] (
	.clk(clk),
	.d(\Add3~80_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[2]~q ),
	.prn(vcc));
defparam \stage_counter[2] .is_wysiwyg = "true";
defparam \stage_counter[2] .power_up = "low";

cycloneiii_lcell_comb \Add3~83 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_refresh_done~q ),
	.datac(\ac_state.s_0~q ),
	.datad(\state.s_dummy_wait~q ),
	.cin(gnd),
	.combout(\Add3~83_combout ),
	.cout());
defparam \Add3~83 .lut_mask = 16'hFFFE;
defparam \Add3~83 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~84 (
	.dataa(\stage_counter[17]~121_combout ),
	.datab(\Add3~83_combout ),
	.datac(\ac_state.s_1~q ),
	.datad(\Add3~61_combout ),
	.cin(gnd),
	.combout(\Add3~84_combout ),
	.cout());
defparam \Add3~84 .lut_mask = 16'hEFFF;
defparam \Add3~84 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add3~85 (
	.dataa(\Add3~82_combout ),
	.datab(\stage_counter[1]~q ),
	.datac(\Add3~60_combout ),
	.datad(\Add3~84_combout ),
	.cin(gnd),
	.combout(\Add3~85_combout ),
	.cout());
defparam \Add3~85 .lut_mask = 16'hFFFE;
defparam \Add3~85 .sum_lutc_input = "datac";

dffeas \stage_counter[1] (
	.clk(clk),
	.d(\Add3~85_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[1]~q ),
	.prn(vcc));
defparam \stage_counter[1] .is_wysiwyg = "true";
defparam \stage_counter[1] .power_up = "low";

cycloneiii_lcell_comb \stage_counter_zero~5 (
	.dataa(gnd),
	.datab(\stage_counter[3]~q ),
	.datac(\stage_counter[2]~q ),
	.datad(\stage_counter[1]~q ),
	.cin(gnd),
	.combout(\stage_counter_zero~5_combout ),
	.cout());
defparam \stage_counter_zero~5 .lut_mask = 16'h3FFF;
defparam \stage_counter_zero~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \stage_counter_zero~6 (
	.dataa(\stage_counter_zero~2_combout ),
	.datab(\stage_counter_zero~3_combout ),
	.datac(\stage_counter_zero~4_combout ),
	.datad(\stage_counter_zero~5_combout ),
	.cin(gnd),
	.combout(\stage_counter_zero~6_combout ),
	.cout());
defparam \stage_counter_zero~6 .lut_mask = 16'h7FFF;
defparam \stage_counter_zero~6 .sum_lutc_input = "datac";

dffeas stage_counter_zero(
	.clk(clk),
	.d(\stage_counter_zero~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter_zero~q ),
	.prn(vcc));
defparam stage_counter_zero.is_wysiwyg = "true";
defparam stage_counter_zero.power_up = "low";

cycloneiii_lcell_comb \process_12~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\process_12~2_combout ),
	.cout());
defparam \process_12~2 .lut_mask = 16'h0FFF;
defparam \process_12~2 .sum_lutc_input = "datac";

dffeas \per_cs_init_seen[0] (
	.clk(clk),
	.d(\Selector216~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_12~2_combout ),
	.q(\per_cs_init_seen[0]~q ),
	.prn(vcc));
defparam \per_cs_init_seen[0] .is_wysiwyg = "true";
defparam \per_cs_init_seen[0] .power_up = "low";

dffeas mem_init_complete(
	.clk(clk),
	.d(\per_cs_init_seen[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_init_complete~q ),
	.prn(vcc));
defparam mem_init_complete.is_wysiwyg = "true";
defparam mem_init_complete.power_up = "low";

cycloneiii_lcell_comb \Selector4~1 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\mem_init_complete~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFEFE;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~2 (
	.dataa(\Selector4~0_combout ),
	.datab(\finished_state~q ),
	.datac(\Selector4~1_combout ),
	.datad(\refreshes_maxed~q ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
defparam \Selector4~2 .lut_mask = 16'hFEFF;
defparam \Selector4~2 .sum_lutc_input = "datac";

dffeas \state.s_topup_refresh (
	.clk(clk),
	.d(\Selector4~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_topup_refresh~q ),
	.prn(vcc));
defparam \state.s_topup_refresh .is_wysiwyg = "true";
defparam \state.s_topup_refresh .power_up = "low";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\state.s_topup_refresh~q ),
	.datac(\finished_state~q ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hFFAC;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \state.s_topup_refresh_done (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_topup_refresh_done~q ),
	.prn(vcc));
defparam \state.s_topup_refresh_done .is_wysiwyg = "true";
defparam \state.s_topup_refresh_done .power_up = "low";

cycloneiii_lcell_comb \refresh_done~2 (
	.dataa(\ac_state.s_0~q ),
	.datab(\state.s_topup_refresh_done~q ),
	.datac(\state.s_refresh_done~q ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\refresh_done~2_combout ),
	.cout());
defparam \refresh_done~2 .lut_mask = 16'hFFFD;
defparam \refresh_done~2 .sum_lutc_input = "datac";

dffeas refresh_done(
	.clk(clk),
	.d(\refresh_done~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_done~q ),
	.prn(vcc));
defparam refresh_done.is_wysiwyg = "true";
defparam refresh_done.power_up = "low";

cycloneiii_lcell_comb \num_stacked_refreshes~9 (
	.dataa(\refresh_due~q ),
	.datab(\num_stacked_refreshes[1]~q ),
	.datac(\num_stacked_refreshes[0]~q ),
	.datad(\refresh_done~q ),
	.cin(gnd),
	.combout(\num_stacked_refreshes~9_combout ),
	.cout());
defparam \num_stacked_refreshes~9 .lut_mask = 16'hFFFE;
defparam \num_stacked_refreshes~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \num_stacked_refreshes~10 (
	.dataa(ctl_init_success),
	.datab(\num_stacked_refreshes[2]~q ),
	.datac(\refresh_due~q ),
	.datad(\num_stacked_refreshes~9_combout ),
	.cin(gnd),
	.combout(\num_stacked_refreshes~10_combout ),
	.cout());
defparam \num_stacked_refreshes~10 .lut_mask = 16'hFFDF;
defparam \num_stacked_refreshes~10 .sum_lutc_input = "datac";

dffeas \num_stacked_refreshes[2] (
	.clk(clk),
	.d(\num_stacked_refreshes~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[2]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[2] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[2] .power_up = "low";

cycloneiii_lcell_comb \LessThan0~0 (
	.dataa(gnd),
	.datab(\num_stacked_refreshes[2]~q ),
	.datac(\num_stacked_refreshes[1]~q ),
	.datad(\num_stacked_refreshes[0]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFC;
defparam \LessThan0~0 .sum_lutc_input = "datac";

dffeas refreshes_maxed(
	.clk(clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refreshes_maxed~q ),
	.prn(vcc));
defparam refreshes_maxed.is_wysiwyg = "true";
defparam refreshes_maxed.power_up = "low";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(\state.s_topup_refresh_done~q ),
	.datab(\finished_state~q ),
	.datac(\refreshes_maxed~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFEFE;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~2 (
	.dataa(dgwb_ac_access_req),
	.datab(dgrb_ac_access_req),
	.datac(curr_cmdcmd_prep_customer_mr_setup),
	.datad(\admin_req_extended~q ),
	.cin(gnd),
	.combout(\Selector7~2_combout ),
	.cout());
defparam \Selector7~2 .lut_mask = 16'h6FFF;
defparam \Selector7~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~3 (
	.dataa(\state.s_access_act~q ),
	.datab(\Selector7~0_combout ),
	.datac(\Selector7~2_combout ),
	.datad(\Selector7~1_combout ),
	.cin(gnd),
	.combout(\Selector7~3_combout ),
	.cout());
defparam \Selector7~3 .lut_mask = 16'hFFFE;
defparam \Selector7~3 .sum_lutc_input = "datac";

dffeas \state.s_access_act (
	.clk(clk),
	.d(\Selector7~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access_act~q ),
	.prn(vcc));
defparam \state.s_access_act .is_wysiwyg = "true";
defparam \state.s_access_act .power_up = "low";

cycloneiii_lcell_comb \WideOr43~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_access_act~q ),
	.datad(\state.s_access_precharge~q ),
	.cin(gnd),
	.combout(\WideOr43~0_combout ),
	.cout());
defparam \WideOr43~0 .lut_mask = 16'h0FFF;
defparam \WideOr43~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector219~7 (
	.dataa(\state.s_topup_refresh~q ),
	.datab(\state.s_refresh~q ),
	.datac(\WideOr41~0_combout ),
	.datad(\WideOr43~0_combout ),
	.cin(gnd),
	.combout(\Selector219~7_combout ),
	.cout());
defparam \Selector219~7 .lut_mask = 16'hEFFF;
defparam \Selector219~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector219~6 (
	.dataa(\ac_state.s_1~q ),
	.datab(\Selector219~7_combout ),
	.datac(\ac_state.s_2~q ),
	.datad(\state~166_combout ),
	.cin(gnd),
	.combout(\Selector219~6_combout ),
	.cout());
defparam \Selector219~6 .lut_mask = 16'hFEFF;
defparam \Selector219~6 .sum_lutc_input = "datac";

dffeas \ac_state.s_2 (
	.clk(clk),
	.d(\Selector219~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_12~2_combout ),
	.q(\ac_state.s_2~q ),
	.prn(vcc));
defparam \ac_state.s_2 .is_wysiwyg = "true";
defparam \ac_state.s_2 .power_up = "low";

cycloneiii_lcell_comb \addr_cmd~507 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.s_topup_refresh~q ),
	.datad(\state.s_refresh~q ),
	.cin(gnd),
	.combout(\addr_cmd~507_combout ),
	.cout());
defparam \addr_cmd~507 .lut_mask = 16'h0FFF;
defparam \addr_cmd~507 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \finished_state~3 (
	.dataa(\finished_state~2_combout ),
	.datab(\ac_state.s_2~q ),
	.datac(\addr_cmd~507_combout ),
	.datad(\WideOr43~0_combout ),
	.cin(gnd),
	.combout(\finished_state~3_combout ),
	.cout());
defparam \finished_state~3 .lut_mask = 16'hEFFF;
defparam \finished_state~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \finished_state~4 (
	.dataa(\process_12~2_combout ),
	.datab(\finished_state~3_combout ),
	.datac(\ac_state.s_7~q ),
	.datad(\state.s_prog_user_mrs~q ),
	.cin(gnd),
	.combout(\finished_state~4_combout ),
	.cout());
defparam \finished_state~4 .lut_mask = 16'hFFFE;
defparam \finished_state~4 .sum_lutc_input = "datac";

dffeas finished_state(
	.clk(clk),
	.d(\finished_state~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_state~q ),
	.prn(vcc));
defparam finished_state.is_wysiwyg = "true";
defparam finished_state.power_up = "low";

cycloneiii_lcell_comb \Selector13~0 (
	.dataa(\state.s_refresh_done~q ),
	.datab(\state.s_refresh~q ),
	.datac(\finished_state~q ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hFFAC;
defparam \Selector13~0 .sum_lutc_input = "datac";

dffeas \state.s_refresh_done (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_refresh_done~q ),
	.prn(vcc));
defparam \state.s_refresh_done .is_wysiwyg = "true";
defparam \state.s_refresh_done .power_up = "low";

cycloneiii_lcell_comb \Selector12~0 (
	.dataa(\state.s_dummy_wait~q ),
	.datab(\state.s_refresh_done~q ),
	.datac(gnd),
	.datad(\refreshes_maxed~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hEEFF;
defparam \Selector12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~1 (
	.dataa(\state.s_refresh~q ),
	.datab(\Selector12~0_combout ),
	.datac(\finished_state~q ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
defparam \Selector12~1 .lut_mask = 16'hFFAC;
defparam \Selector12~1 .sum_lutc_input = "datac";

dffeas \state.s_refresh (
	.clk(clk),
	.d(\Selector12~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(ctl_init_success),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_refresh~q ),
	.prn(vcc));
defparam \state.s_refresh .is_wysiwyg = "true";
defparam \state.s_refresh .power_up = "low";

cycloneiii_lcell_comb WideOr45(
	.dataa(\state.s_dummy_wait~q ),
	.datab(\state.s_topup_refresh_done~q ),
	.datac(\state.s_refresh_done~q ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\WideOr45~combout ),
	.cout());
defparam WideOr45.lut_mask = 16'hFEFF;
defparam WideOr45.sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector286~5 (
	.dataa(\state.s_topup_refresh~q ),
	.datab(\state.s_refresh~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\WideOr45~combout ),
	.cin(gnd),
	.combout(\Selector286~5_combout ),
	.cout());
defparam \Selector286~5 .lut_mask = 16'hF7FF;
defparam \Selector286~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector286~4 (
	.dataa(\addr_cmd[0].cke[0]~0_combout ),
	.datab(\Selector286~2_combout ),
	.datac(\Selector286~5_combout ),
	.datad(\Selector286~3_combout ),
	.cin(gnd),
	.combout(\Selector286~4_combout ),
	.cout());
defparam \Selector286~4 .lut_mask = 16'hFFFE;
defparam \Selector286~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector302~3 (
	.dataa(addr_cmd0cs_n0),
	.datab(\state.s_run_init_seq~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector302~3_combout ),
	.cout());
defparam \Selector302~3 .lut_mask = 16'hEEEE;
defparam \Selector302~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~508 (
	.dataa(\addr_cmd~507_combout ),
	.datab(\ac_state.s_1~q ),
	.datac(\WideOr45~combout ),
	.datad(\Selector302~3_combout ),
	.cin(gnd),
	.combout(\addr_cmd~508_combout ),
	.cout());
defparam \addr_cmd~508 .lut_mask = 16'hBFFF;
defparam \addr_cmd~508 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector302~4 (
	.dataa(addr_cmd0cs_n0),
	.datab(\state.s_run_init_seq~q ),
	.datac(\ac_state.s_1~q ),
	.datad(\state.s_access_act~q ),
	.cin(gnd),
	.combout(\Selector302~4_combout ),
	.cout());
defparam \Selector302~4 .lut_mask = 16'h7FFF;
defparam \Selector302~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~1 (
	.dataa(\state.s_access_precharge~q ),
	.datab(\ac_state.s_1~q ),
	.datac(\ac_state.s_0~q ),
	.datad(\ac_state.s_2~q ),
	.cin(gnd),
	.combout(\Selector269~1_combout ),
	.cout());
defparam \Selector269~1 .lut_mask = 16'hEFFF;
defparam \Selector269~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~509 (
	.dataa(\Selector302~5_combout ),
	.datab(\Selector302~4_combout ),
	.datac(\ac_state.s_0~q ),
	.datad(\Selector269~1_combout ),
	.cin(gnd),
	.combout(\addr_cmd~509_combout ),
	.cout());
defparam \addr_cmd~509 .lut_mask = 16'hEFFF;
defparam \addr_cmd~509 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~510 (
	.dataa(\Selector302~2_combout ),
	.datab(\addr_cmd~508_combout ),
	.datac(\addr_cmd~509_combout ),
	.datad(\process_12~2_combout ),
	.cin(gnd),
	.combout(\addr_cmd~510_combout ),
	.cout());
defparam \addr_cmd~510 .lut_mask = 16'hFFFE;
defparam \addr_cmd~510 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_10~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\WideNor0~0_combout ),
	.cout());
defparam \WideNor0~0 .lut_mask = 16'h0FFF;
defparam \WideNor0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~511 (
	.dataa(\addr_cmd~510_combout ),
	.datab(\process_12~2_combout ),
	.datac(\WideNor0~0_combout ),
	.datad(\Selector302~3_combout ),
	.cin(gnd),
	.combout(\addr_cmd~511_combout ),
	.cout());
defparam \addr_cmd~511 .lut_mask = 16'hFFFD;
defparam \addr_cmd~511 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~512 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(\state.s_access_precharge~q ),
	.datac(gnd),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\addr_cmd~512_combout ),
	.cout());
defparam \addr_cmd~512 .lut_mask = 16'hEEFF;
defparam \addr_cmd~512 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~2 (
	.dataa(\state.s_run_init_seq~q ),
	.datab(\ac_state.s_10~q ),
	.datac(\process_12~6_combout ),
	.datad(\state.s_reset~q ),
	.cin(gnd),
	.combout(\Selector269~2_combout ),
	.cout());
defparam \Selector269~2 .lut_mask = 16'hFFFE;
defparam \Selector269~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~0 (
	.dataa(\ac_state.s_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_state.s_8~q ),
	.cin(gnd),
	.combout(\Selector269~0_combout ),
	.cout());
defparam \Selector269~0 .lut_mask = 16'hAAFF;
defparam \Selector269~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~551 (
	.dataa(\ac_state.s_6~q ),
	.datab(\ac_state.s_5~q ),
	.datac(\state.s_program_cal_mrs~q ),
	.datad(\Selector269~0_combout ),
	.cin(gnd),
	.combout(\addr_cmd~551_combout ),
	.cout());
defparam \addr_cmd~551 .lut_mask = 16'hFEFF;
defparam \addr_cmd~551 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~514 (
	.dataa(\addr_cmd~513_combout ),
	.datab(\state.s_access~q ),
	.datac(\addr_cmd~551_combout ),
	.datad(\state.s_idle~q ),
	.cin(gnd),
	.combout(\addr_cmd~514_combout ),
	.cout());
defparam \addr_cmd~514 .lut_mask = 16'hBFFF;
defparam \addr_cmd~514 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~515 (
	.dataa(\process_12~2_combout ),
	.datab(\addr_cmd~512_combout ),
	.datac(\Selector269~2_combout ),
	.datad(\addr_cmd~514_combout ),
	.cin(gnd),
	.combout(\addr_cmd~515_combout ),
	.cout());
defparam \addr_cmd~515 .lut_mask = 16'hFEFF;
defparam \addr_cmd~515 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~215 (
	.dataa(\ac_state.s_2~q ),
	.datab(\ac_state.s_0~q ),
	.datac(gnd),
	.datad(\ac_state.s_1~q ),
	.cin(gnd),
	.combout(\addr_cmd~215_combout ),
	.cout());
defparam \addr_cmd~215 .lut_mask = 16'hEEFF;
defparam \addr_cmd~215 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~516 (
	.dataa(\WideOr32~0_combout ),
	.datab(\WideOr26~combout ),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\WideOr45~combout ),
	.cin(gnd),
	.combout(\addr_cmd~516_combout ),
	.cout());
defparam \addr_cmd~516 .lut_mask = 16'hBFFF;
defparam \addr_cmd~516 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~517 (
	.dataa(\process_12~2_combout ),
	.datab(\addr_cmd~516_combout ),
	.datac(\WideOr26~0_combout ),
	.datad(\state.s_program_cal_mrs~q ),
	.cin(gnd),
	.combout(\addr_cmd~517_combout ),
	.cout());
defparam \addr_cmd~517 .lut_mask = 16'hFEFF;
defparam \addr_cmd~517 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~518 (
	.dataa(\state.s_reset~q ),
	.datab(\state.s_access_precharge~q ),
	.datac(\addr_cmd~215_combout ),
	.datad(\addr_cmd~517_combout ),
	.cin(gnd),
	.combout(\addr_cmd~518_combout ),
	.cout());
defparam \addr_cmd~518 .lut_mask = 16'hFEFF;
defparam \addr_cmd~518 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~519 (
	.dataa(addr_cmd0addr0),
	.datab(\addr_cmd~515_combout ),
	.datac(\addr_cmd~518_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr_cmd~519_combout ),
	.cout());
defparam \addr_cmd~519 .lut_mask = 16'hFEFE;
defparam \addr_cmd~519 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~520 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(gnd),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~520_combout ),
	.cout());
defparam \addr_cmd~520 .lut_mask = 16'hAFFF;
defparam \addr_cmd~520 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~521 (
	.dataa(\ac_state.s_5~q ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~521_combout ),
	.cout());
defparam \addr_cmd~521 .lut_mask = 16'hEFFF;
defparam \addr_cmd~521 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~522 (
	.dataa(\ac_state.s_3~q ),
	.datab(\ac_state.s_7~q ),
	.datac(\addr_cmd~520_combout ),
	.datad(\addr_cmd~521_combout ),
	.cin(gnd),
	.combout(\addr_cmd~522_combout ),
	.cout());
defparam \addr_cmd~522 .lut_mask = 16'h7FFF;
defparam \addr_cmd~522 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~523 (
	.dataa(addr_cmd0addr1),
	.datab(\addr_cmd~515_combout ),
	.datac(\addr_cmd~518_combout ),
	.datad(\addr_cmd~522_combout ),
	.cin(gnd),
	.combout(\addr_cmd~523_combout ),
	.cout());
defparam \addr_cmd~523 .lut_mask = 16'hFEFF;
defparam \addr_cmd~523 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~524 (
	.dataa(addr_cmd0addr4),
	.datab(\addr_cmd~515_combout ),
	.datac(\addr_cmd~518_combout ),
	.datad(\addr_cmd~522_combout ),
	.cin(gnd),
	.combout(\addr_cmd~524_combout ),
	.cout());
defparam \addr_cmd~524 .lut_mask = 16'hFEFF;
defparam \addr_cmd~524 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~525 (
	.dataa(\ac_state.s_3~q ),
	.datab(\state.s_program_cal_mrs~q ),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~525_combout ),
	.cout());
defparam \addr_cmd~525 .lut_mask = 16'hEFFF;
defparam \addr_cmd~525 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~526 (
	.dataa(\addr_cmd~525_combout ),
	.datab(addr_cmd0addr8),
	.datac(\addr_cmd~515_combout ),
	.datad(\addr_cmd~518_combout ),
	.cin(gnd),
	.combout(\addr_cmd~526_combout ),
	.cout());
defparam \addr_cmd~526 .lut_mask = 16'hFFFE;
defparam \addr_cmd~526 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~527 (
	.dataa(addr_cmd0addr10),
	.datab(\state.s_reset~q ),
	.datac(\state.s_access_precharge~q ),
	.datad(\addr_cmd~517_combout ),
	.cin(gnd),
	.combout(\addr_cmd~527_combout ),
	.cout());
defparam \addr_cmd~527 .lut_mask = 16'hFEFF;
defparam \addr_cmd~527 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_state~96 (
	.dataa(\ac_state.s_2~q ),
	.datab(\ac_state~93_combout ),
	.datac(\state.s_run_init_seq~q ),
	.datad(\process_12~6_combout ),
	.cin(gnd),
	.combout(\ac_state~96_combout ),
	.cout());
defparam \ac_state~96 .lut_mask = 16'hFFFE;
defparam \ac_state~96 .sum_lutc_input = "datac";

dffeas \ac_state.s_3 (
	.clk(clk),
	.d(\ac_state~96_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_state~91_combout ),
	.q(\ac_state.s_3~q ),
	.prn(vcc));
defparam \ac_state.s_3 .is_wysiwyg = "true";
defparam \ac_state.s_3 .power_up = "low";

cycloneiii_lcell_comb \Selector221~1 (
	.dataa(\Selector221~0_combout ),
	.datab(\ac_state.s_3~q ),
	.datac(\state.s_prog_user_mrs~q ),
	.datad(\WideOr41~0_combout ),
	.cin(gnd),
	.combout(\Selector221~1_combout ),
	.cout());
defparam \Selector221~1 .lut_mask = 16'hFEFF;
defparam \Selector221~1 .sum_lutc_input = "datac";

dffeas \ac_state.s_4 (
	.clk(clk),
	.d(\Selector221~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_12~2_combout ),
	.q(\ac_state.s_4~q ),
	.prn(vcc));
defparam \ac_state.s_4 .is_wysiwyg = "true";
defparam \ac_state.s_4 .power_up = "low";

cycloneiii_lcell_comb \addr_cmd~528 (
	.dataa(\Selector269~2_combout ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\ac_state.s_0~q ),
	.datad(\addr_cmd~514_combout ),
	.cin(gnd),
	.combout(\addr_cmd~528_combout ),
	.cout());
defparam \addr_cmd~528 .lut_mask = 16'hEFFF;
defparam \addr_cmd~528 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~529 (
	.dataa(\Selector269~1_combout ),
	.datab(addr_cmd0addr10),
	.datac(\ac_state.s_0~q ),
	.datad(\addr_cmd~528_combout ),
	.cin(gnd),
	.combout(\addr_cmd~529_combout ),
	.cout());
defparam \addr_cmd~529 .lut_mask = 16'hFFFE;
defparam \addr_cmd~529 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~530 (
	.dataa(\process_12~2_combout ),
	.datab(\ac_state.s_1~q ),
	.datac(\stage_counter[17]~118_combout ),
	.datad(\addr_cmd~529_combout ),
	.cin(gnd),
	.combout(\addr_cmd~530_combout ),
	.cout());
defparam \addr_cmd~530 .lut_mask = 16'hFFFE;
defparam \addr_cmd~530 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~531 (
	.dataa(\addr_cmd~527_combout ),
	.datab(\ac_state.s_4~q ),
	.datac(\addr_cmd~520_combout ),
	.datad(\addr_cmd~530_combout ),
	.cin(gnd),
	.combout(\addr_cmd~531_combout ),
	.cout());
defparam \addr_cmd~531 .lut_mask = 16'hFFFE;
defparam \addr_cmd~531 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~532 (
	.dataa(\state.s_prog_user_mrs~q ),
	.datab(gnd),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~532_combout ),
	.cout());
defparam \addr_cmd~532 .lut_mask = 16'hAFFF;
defparam \addr_cmd~532 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~533 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_3~q ),
	.datad(\ac_state.s_4~q ),
	.cin(gnd),
	.combout(\addr_cmd~533_combout ),
	.cout());
defparam \addr_cmd~533 .lut_mask = 16'h0FFF;
defparam \addr_cmd~533 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~534 (
	.dataa(\ac_state.s_2~q ),
	.datab(\addr_cmd~520_combout ),
	.datac(\addr_cmd~532_combout ),
	.datad(\addr_cmd~533_combout ),
	.cin(gnd),
	.combout(\addr_cmd~534_combout ),
	.cout());
defparam \addr_cmd~534 .lut_mask = 16'hFEFF;
defparam \addr_cmd~534 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~535 (
	.dataa(\addr_cmd~534_combout ),
	.datab(addr_cmd0ba0),
	.datac(\addr_cmd~515_combout ),
	.datad(\addr_cmd~518_combout ),
	.cin(gnd),
	.combout(\addr_cmd~535_combout ),
	.cout());
defparam \addr_cmd~535 .lut_mask = 16'hFFFE;
defparam \addr_cmd~535 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~536 (
	.dataa(\addr_cmd~532_combout ),
	.datab(\ac_state.s_3~q ),
	.datac(\ac_state.s_2~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr_cmd~536_combout ),
	.cout());
defparam \addr_cmd~536 .lut_mask = 16'hFEFE;
defparam \addr_cmd~536 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~537 (
	.dataa(\addr_cmd~536_combout ),
	.datab(addr_cmd0ba1),
	.datac(\addr_cmd~515_combout ),
	.datad(\addr_cmd~518_combout ),
	.cin(gnd),
	.combout(\addr_cmd~537_combout ),
	.cout());
defparam \addr_cmd~537 .lut_mask = 16'hFFFE;
defparam \addr_cmd~537 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector269~9 (
	.dataa(\Selector269~8_combout ),
	.datab(addr_cmd0ras_n),
	.datac(\Selector269~2_combout ),
	.datad(\WideOr38~1_combout ),
	.cin(gnd),
	.combout(\Selector269~9_combout ),
	.cout());
defparam \Selector269~9 .lut_mask = 16'hFEFF;
defparam \Selector269~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~538 (
	.dataa(addr_cmd0ras_n),
	.datab(\Selector269~9_combout ),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~538_combout ),
	.cout());
defparam \addr_cmd~538 .lut_mask = 16'hEFFE;
defparam \addr_cmd~538 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr32~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_state.s_7~q ),
	.datad(\ac_state.s_6~q ),
	.cin(gnd),
	.combout(\WideOr32~0_combout ),
	.cout());
defparam \WideOr32~0 .lut_mask = 16'h0FFF;
defparam \WideOr32~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~543 (
	.dataa(\state.s_program_cal_mrs~q ),
	.datab(addr_cmd0cas_n),
	.datac(\ac_state.s_8~q ),
	.datad(\WideOr32~0_combout ),
	.cin(gnd),
	.combout(\addr_cmd~543_combout ),
	.cout());
defparam \addr_cmd~543 .lut_mask = 16'hFEFF;
defparam \addr_cmd~543 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~540 (
	.dataa(addr_cmd0cas_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\addr_cmd~540_combout ),
	.cout());
defparam \addr_cmd~540 .lut_mask = 16'hAAFF;
defparam \addr_cmd~540 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~544 (
	.dataa(\state.s_access_precharge~q ),
	.datab(\addr_cmd~540_combout ),
	.datac(\ac_state.s_1~q ),
	.datad(\addr_cmd~507_combout ),
	.cin(gnd),
	.combout(\addr_cmd~544_combout ),
	.cout());
defparam \addr_cmd~544 .lut_mask = 16'hFEFF;
defparam \addr_cmd~544 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~545 (
	.dataa(\ac_state.s_4~q ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(addr_cmd0cas_n),
	.datad(\WideOr38~1_combout ),
	.cin(gnd),
	.combout(\addr_cmd~545_combout ),
	.cout());
defparam \addr_cmd~545 .lut_mask = 16'hFEFF;
defparam \addr_cmd~545 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~546 (
	.dataa(\addr_cmd~542_combout ),
	.datab(\addr_cmd~543_combout ),
	.datac(\addr_cmd~544_combout ),
	.datad(\addr_cmd~545_combout ),
	.cin(gnd),
	.combout(\addr_cmd~546_combout ),
	.cout());
defparam \addr_cmd~546 .lut_mask = 16'hFFFE;
defparam \addr_cmd~546 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~547 (
	.dataa(\process_12~2_combout ),
	.datab(\addr_cmd~546_combout ),
	.datac(addr_cmd0cas_n),
	.datad(\Selector269~2_combout ),
	.cin(gnd),
	.combout(\addr_cmd~547_combout ),
	.cout());
defparam \addr_cmd~547 .lut_mask = 16'hFFFE;
defparam \addr_cmd~547 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~548 (
	.dataa(\state.s_access_precharge~q ),
	.datab(\addr_cmd~215_combout ),
	.datac(\addr_cmd~507_combout ),
	.datad(\addr_cmd~517_combout ),
	.cin(gnd),
	.combout(\addr_cmd~548_combout ),
	.cout());
defparam \addr_cmd~548 .lut_mask = 16'hEFFF;
defparam \addr_cmd~548 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~549 (
	.dataa(\addr_cmd~547_combout ),
	.datab(addr_cmd0cas_n),
	.datac(\state.s_reset~q ),
	.datad(\addr_cmd~548_combout ),
	.cin(gnd),
	.combout(\addr_cmd~549_combout ),
	.cout());
defparam \addr_cmd~549 .lut_mask = 16'hFFFE;
defparam \addr_cmd~549 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~0 (
	.dataa(\Selector269~1_combout ),
	.datab(\state.s_prog_user_mrs~q ),
	.datac(\WideOr32~0_combout ),
	.datad(\WideOr26~combout ),
	.cin(gnd),
	.combout(\Selector270~0_combout ),
	.cout());
defparam \Selector270~0 .lut_mask = 16'hFEFF;
defparam \Selector270~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~6 (
	.dataa(\Selector270~5_combout ),
	.datab(\Selector270~0_combout ),
	.datac(addr_cmd0we_n),
	.datad(\ac_state.s_0~q ),
	.cin(gnd),
	.combout(\Selector270~6_combout ),
	.cout());
defparam \Selector270~6 .lut_mask = 16'hFFFE;
defparam \Selector270~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector270~7 (
	.dataa(\Selector270~4_combout ),
	.datab(\Selector270~6_combout ),
	.datac(addr_cmd0we_n),
	.datad(\Selector269~2_combout ),
	.cin(gnd),
	.combout(\Selector270~7_combout ),
	.cout());
defparam \Selector270~7 .lut_mask = 16'hFFFE;
defparam \Selector270~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \addr_cmd~550 (
	.dataa(addr_cmd0we_n),
	.datab(\Selector270~7_combout ),
	.datac(\state.s_reset~q ),
	.datad(\stage_counter_zero~q ),
	.cin(gnd),
	.combout(\addr_cmd~550_combout ),
	.cout());
defparam \addr_cmd~550 .lut_mask = 16'hEFFE;
defparam \addr_cmd~550 .sum_lutc_input = "datac";

dffeas command_done(
	.clk(clk),
	.d(\stage_counter[17]~118_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\finished_state~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\command_done~q ),
	.prn(vcc));
defparam command_done.is_wysiwyg = "true";
defparam command_done.power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_ctrl (
	clk,
	rst_n,
	ctl_init_success1,
	states_init_dram,
	WideOr34,
	ac_muxctrl_broadcast_rcommandcmd_init_dram,
	admin_ctrlcommand_done,
	dgwb_ctrlcommand_done,
	curr_cmdcmd_prep_customer_mr_setup,
	Selector1,
	curr_cmdcmd_write_btp,
	curr_cmdcmd_write_mtp,
	curr_cmdcmd_was,
	WideOr0,
	dgrb_ctrlcommand_done,
	curr_cmdcmd_idle,
	WideOr11,
	last_states_rdv,
	last_states_read_mtp,
	last_states_rrp_seek,
	last_states_adv_rd_lat,
	last_states_rrp_sweep,
	last_states_adv_wr_lat,
	last_states_rrp_reset,
	Selector58,
	ctrl_op_reccommand_opsingle_bit,
	ctrl_op_reccommand_opmtp_almt,
	Selector57,
	Selector52,
	dgrb_ctrlcommand_result_5,
	dgrb_ctrlcommand_result_4,
	dgrb_ctrlcommand_result_3,
	dgrb_ctrlcommand_result_2,
	dgrb_ctrlcommand_result_1,
	dgrb_ctrlcommand_result_0,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	rst_n;
output 	ctl_init_success1;
output 	states_init_dram;
output 	WideOr34;
input 	ac_muxctrl_broadcast_rcommandcmd_init_dram;
input 	admin_ctrlcommand_done;
input 	dgwb_ctrlcommand_done;
output 	curr_cmdcmd_prep_customer_mr_setup;
output 	Selector1;
output 	curr_cmdcmd_write_btp;
output 	curr_cmdcmd_write_mtp;
output 	curr_cmdcmd_was;
output 	WideOr0;
input 	dgrb_ctrlcommand_done;
output 	curr_cmdcmd_idle;
output 	WideOr11;
output 	last_states_rdv;
output 	last_states_read_mtp;
output 	last_states_rrp_seek;
output 	last_states_adv_rd_lat;
output 	last_states_rrp_sweep;
output 	last_states_adv_wr_lat;
output 	last_states_rrp_reset;
output 	Selector58;
output 	ctrl_op_reccommand_opsingle_bit;
output 	ctrl_op_reccommand_opmtp_almt;
output 	Selector57;
output 	Selector52;
input 	dgrb_ctrlcommand_result_5;
input 	dgrb_ctrlcommand_result_4;
input 	dgrb_ctrlcommand_result_3;
input 	dgrb_ctrlcommand_result_2;
input 	dgrb_ctrlcommand_result_1;
input 	dgrb_ctrlcommand_result_0;
input 	GND_port;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \dll_lock_counter[1]~q ;
wire \dll_lock_counter[2]~q ;
wire \dll_lock_counter[3]~q ;
wire \dll_lock_counter[4]~q ;
wire \dll_lock_counter[5]~q ;
wire \dll_lock_counter[6]~q ;
wire \dll_lock_counter[7]~q ;
wire \dll_lock_counter[10]~q ;
wire \dll_lock_counter[9]~q ;
wire \dll_lock_counter[8]~q ;
wire \tracking_ms_counter[0]~q ;
wire \tracking_ms_counter[1]~q ;
wire \tracking_ms_counter[4]~q ;
wire \dll_lock_counter[1]~34_cout ;
wire \dll_lock_counter[1]~36 ;
wire \dll_lock_counter[1]~35_combout ;
wire \dll_lock_counter[2]~38 ;
wire \dll_lock_counter[2]~37_combout ;
wire \dll_lock_counter[3]~40 ;
wire \dll_lock_counter[3]~39_combout ;
wire \dll_lock_counter[4]~42 ;
wire \dll_lock_counter[4]~41_combout ;
wire \dll_lock_counter[5]~44 ;
wire \dll_lock_counter[5]~43_combout ;
wire \dll_lock_counter[6]~46 ;
wire \dll_lock_counter[6]~45_combout ;
wire \dll_lock_counter[7]~48 ;
wire \dll_lock_counter[7]~47_combout ;
wire \dll_lock_counter[8]~50 ;
wire \dll_lock_counter[8]~49_combout ;
wire \dll_lock_counter[9]~52 ;
wire \dll_lock_counter[9]~51_combout ;
wire \dll_lock_counter[10]~53_combout ;
wire \tracking_ms_counter[0]~40_combout ;
wire \tracking_ms_counter[1]~44_combout ;
wire \tracking_ms_counter[4]~50_combout ;
wire \Add7~3 ;
wire \Add7~5 ;
wire \Add7~4_combout ;
wire \Add7~7 ;
wire \Add7~6_combout ;
wire \Add7~9 ;
wire \Add7~8_combout ;
wire \Add7~11 ;
wire \Add7~10_combout ;
wire \Add7~13 ;
wire \Add7~12_combout ;
wire \Add7~15 ;
wire \Add7~14_combout ;
wire \Add7~17 ;
wire \Add7~16_combout ;
wire \Add7~19 ;
wire \Add7~18_combout ;
wire \Add7~21 ;
wire \Add7~20_combout ;
wire \Add7~23 ;
wire \Add7~22_combout ;
wire \Add7~25 ;
wire \Add7~24_combout ;
wire \Add7~27 ;
wire \Add7~26_combout ;
wire \Add7~29 ;
wire \Add7~28_combout ;
wire \Add7~31 ;
wire \Add7~30_combout ;
wire \Add7~33 ;
wire \Add7~32_combout ;
wire \Add7~34_combout ;
wire \curr_ctrl.command_done~q ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \dll_lock_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \WideNor1~0_combout ;
wire \WideNor1~1_combout ;
wire \last_state.s_reset~q ;
wire \WideNor1~2_combout ;
wire \last_state.s_cal~q ;
wire \WideNor1~3_combout ;
wire \WideNor1~4_combout ;
wire \WideNor1~5_combout ;
wire \Equal5~0_combout ;
wire \milisecond_tick_gen_count[17]~q ;
wire \milisecond_tick_gen_count[14]~q ;
wire \milisecond_tick_gen_count[16]~q ;
wire \milisecond_tick_gen_count[15]~q ;
wire \Equal4~0_combout ;
wire \milisecond_tick_gen_count[11]~q ;
wire \milisecond_tick_gen_count[13]~q ;
wire \milisecond_tick_gen_count[12]~q ;
wire \milisecond_tick_gen_count[10]~q ;
wire \Equal4~1_combout ;
wire \milisecond_tick_gen_count[8]~q ;
wire \milisecond_tick_gen_count[7]~q ;
wire \milisecond_tick_gen_count[6]~q ;
wire \milisecond_tick_gen_count[9]~q ;
wire \Equal4~2_combout ;
wire \milisecond_tick_gen_count[5]~q ;
wire \milisecond_tick_gen_count[2]~q ;
wire \milisecond_tick_gen_count[4]~q ;
wire \milisecond_tick_gen_count[3]~q ;
wire \Equal4~3_combout ;
wire \Equal4~4_combout ;
wire \WideNor1~12_combout ;
wire \dll_lock_counter[0]~32_combout ;
wire \milisecond_tick_gen_count[17]~74_combout ;
wire \milisecond_tick_gen_count[14]~75_combout ;
wire \milisecond_tick_gen_count[0]~76_combout ;
wire \milisecond_tick_gen_count[16]~77_combout ;
wire \milisecond_tick_gen_count[15]~78_combout ;
wire \milisecond_tick_gen_count[11]~79_combout ;
wire \milisecond_tick_gen_count[13]~80_combout ;
wire \milisecond_tick_gen_count[12]~81_combout ;
wire \milisecond_tick_gen_count[10]~82_combout ;
wire \milisecond_tick_gen_count[8]~83_combout ;
wire \milisecond_tick_gen_count[7]~84_combout ;
wire \milisecond_tick_gen_count[6]~85_combout ;
wire \milisecond_tick_gen_count[9]~86_combout ;
wire \milisecond_tick_gen_count[5]~87_combout ;
wire \milisecond_tick_gen_count[2]~88_combout ;
wire \milisecond_tick_gen_count[4]~89_combout ;
wire \milisecond_tick_gen_count[3]~90_combout ;
wire \mtp_almt:dvw_size_a0[5]~q ;
wire \mtp_almt:dvw_size_a0[4]~q ;
wire \mtp_almt:dvw_size_a0[3]~q ;
wire \mtp_almt:dvw_size_a0[2]~q ;
wire \mtp_almt:dvw_size_a0[1]~q ;
wire \mtp_almt:dvw_size_a0[0]~q ;
wire \mtp_almt:dvw_size_a0[0]~0_combout ;
wire \tracking_ms_counter[0]~41 ;
wire \tracking_ms_counter[1]~45 ;
wire \tracking_ms_counter[2]~47 ;
wire \tracking_ms_counter[3]~49 ;
wire \tracking_ms_counter[4]~51 ;
wire \tracking_ms_counter[5]~52_combout ;
wire \Selector34~0_combout ;
wire \last_state.s_tracking~q ;
wire \WideNor1~6_combout ;
wire \state.s_write_btp~q ;
wire \WideNor1~7_combout ;
wire \state~163_combout ;
wire \hold_state~2_combout ;
wire \state.s_read_mtp~q ;
wire \state~46_combout ;
wire \state.s_rrp_reset~q ;
wire \state.s_rrp_sweep~q ;
wire \WideNor1~8_combout ;
wire \WideNor1~9_combout ;
wire \last_state.s_poa~q ;
wire \WideNor1~10_combout ;
wire \process_14~13_combout ;
wire \WideNor1~11_combout ;
wire \WideOr28~0_combout ;
wire \dis_state~5_combout ;
wire \master_ctrl_op_rec~41_combout ;
wire \state.s_phy_initialise~1_combout ;
wire \state.s_phy_initialise~q ;
wire \dis_state~6_combout ;
wire \dis_state~q ;
wire \hold_state~q ;
wire \state~162_combout ;
wire \state.s_cal~q ;
wire \mtp_almts_checked[1]~8_combout ;
wire \mtp_almts_checked[0]~q ;
wire \Selector33~0_combout ;
wire \mtp_almts_checked[1]~q ;
wire \state~164_combout ;
wire \state.s_rrp_seek~q ;
wire \state.s_rdv~q ;
wire \state.s_was~q ;
wire \state.s_adv_rd_lat~q ;
wire \state.s_adv_wr_lat~q ;
wire \state.s_poa~q ;
wire \state.s_tracking_setup~q ;
wire \state.s_prep_customer_mr_setup~q ;
wire \Selector30~0_combout ;
wire \state.s_operational~q ;
wire \last_state.s_operational~q ;
wire \process_16~0_combout ;
wire \milisecond_tick_gen_count[0]~73_combout ;
wire \milisecond_tick_gen_count[0]~92_combout ;
wire \milisecond_tick_gen_count[0]~q ;
wire \Equal4~5_combout ;
wire \milisecond_tick_gen_count[2]~72_combout ;
wire \Add7~1_cout ;
wire \Add7~2_combout ;
wire \milisecond_tick_gen_count[1]~91_combout ;
wire \milisecond_tick_gen_count[1]~q ;
wire \tracking_ms_counter[0]~42_combout ;
wire \tracking_ms_counter[0]~43_combout ;
wire \tracking_ms_counter[5]~q ;
wire \tracking_ms_counter[5]~53 ;
wire \tracking_ms_counter[6]~54_combout ;
wire \tracking_ms_counter[6]~q ;
wire \tracking_ms_counter[6]~55 ;
wire \tracking_ms_counter[7]~56_combout ;
wire \tracking_ms_counter[7]~q ;
wire \Equal5~1_combout ;
wire \tracking_ms_counter[2]~46_combout ;
wire \tracking_ms_counter[2]~q ;
wire \tracking_ms_counter[3]~48_combout ;
wire \tracking_ms_counter[3]~q ;
wire \Equal5~2_combout ;
wire \tracking_update_due~5_combout ;
wire \tracking_update_due~q ;
wire \Selector29~0_combout ;
wire \state.s_tracking~q ;
wire \Selector37~0_combout ;
wire \int_ctl_init_success~q ;
wire \state.s_reset~q ;
wire \WideOr34~6_combout ;
wire \state.s_write_mtp~q ;
wire \WideOr34~7_combout ;
wire \last_state.s_tracking_setup~q ;
wire \last_state.s_phy_initialise~q ;
wire \WideNor1~13_combout ;
wire \WideNor1~14_combout ;
wire \WideNor1~15_combout ;
wire \WideOr1~8_combout ;
wire \WideNor1~16_combout ;
wire \Selector41~0_combout ;
wire \Selector4~0_combout ;
wire \curr_ctrl.command_result[5]~q ;
wire \mtp_almt:dvw_size_a1[0]~0_combout ;
wire \mtp_almt:dvw_size_a1[5]~q ;
wire \Selector5~0_combout ;
wire \curr_ctrl.command_result[4]~q ;
wire \mtp_almt:dvw_size_a1[4]~q ;
wire \Selector6~0_combout ;
wire \curr_ctrl.command_result[3]~q ;
wire \mtp_almt:dvw_size_a1[3]~q ;
wire \Selector7~0_combout ;
wire \curr_ctrl.command_result[2]~q ;
wire \mtp_almt:dvw_size_a1[2]~q ;
wire \Selector8~0_combout ;
wire \curr_ctrl.command_result[1]~q ;
wire \mtp_almt:dvw_size_a1[1]~q ;
wire \Selector9~0_combout ;
wire \curr_ctrl.command_result[0]~q ;
wire \mtp_almt:dvw_size_a1[0]~q ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~10_combout ;
wire \mtp_correct_almt~q ;


dffeas \dll_lock_counter[1] (
	.clk(clk),
	.d(\dll_lock_counter[1]~35_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[1]~q ),
	.prn(vcc));
defparam \dll_lock_counter[1] .is_wysiwyg = "true";
defparam \dll_lock_counter[1] .power_up = "low";

dffeas \dll_lock_counter[2] (
	.clk(clk),
	.d(\dll_lock_counter[2]~37_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[2]~q ),
	.prn(vcc));
defparam \dll_lock_counter[2] .is_wysiwyg = "true";
defparam \dll_lock_counter[2] .power_up = "low";

dffeas \dll_lock_counter[3] (
	.clk(clk),
	.d(\dll_lock_counter[3]~39_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[3]~q ),
	.prn(vcc));
defparam \dll_lock_counter[3] .is_wysiwyg = "true";
defparam \dll_lock_counter[3] .power_up = "low";

dffeas \dll_lock_counter[4] (
	.clk(clk),
	.d(\dll_lock_counter[4]~41_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[4]~q ),
	.prn(vcc));
defparam \dll_lock_counter[4] .is_wysiwyg = "true";
defparam \dll_lock_counter[4] .power_up = "low";

dffeas \dll_lock_counter[5] (
	.clk(clk),
	.d(\dll_lock_counter[5]~43_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[5]~q ),
	.prn(vcc));
defparam \dll_lock_counter[5] .is_wysiwyg = "true";
defparam \dll_lock_counter[5] .power_up = "low";

dffeas \dll_lock_counter[6] (
	.clk(clk),
	.d(\dll_lock_counter[6]~45_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[6]~q ),
	.prn(vcc));
defparam \dll_lock_counter[6] .is_wysiwyg = "true";
defparam \dll_lock_counter[6] .power_up = "low";

dffeas \dll_lock_counter[7] (
	.clk(clk),
	.d(\dll_lock_counter[7]~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[7]~q ),
	.prn(vcc));
defparam \dll_lock_counter[7] .is_wysiwyg = "true";
defparam \dll_lock_counter[7] .power_up = "low";

dffeas \dll_lock_counter[10] (
	.clk(clk),
	.d(\dll_lock_counter[10]~53_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[10]~q ),
	.prn(vcc));
defparam \dll_lock_counter[10] .is_wysiwyg = "true";
defparam \dll_lock_counter[10] .power_up = "low";

dffeas \dll_lock_counter[9] (
	.clk(clk),
	.d(\dll_lock_counter[9]~51_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[9]~q ),
	.prn(vcc));
defparam \dll_lock_counter[9] .is_wysiwyg = "true";
defparam \dll_lock_counter[9] .power_up = "low";

dffeas \dll_lock_counter[8] (
	.clk(clk),
	.d(\dll_lock_counter[8]~49_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~3_combout ),
	.q(\dll_lock_counter[8]~q ),
	.prn(vcc));
defparam \dll_lock_counter[8] .is_wysiwyg = "true";
defparam \dll_lock_counter[8] .power_up = "low";

dffeas \tracking_ms_counter[0] (
	.clk(clk),
	.d(\tracking_ms_counter[0]~40_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[0]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[0] .is_wysiwyg = "true";
defparam \tracking_ms_counter[0] .power_up = "low";

dffeas \tracking_ms_counter[1] (
	.clk(clk),
	.d(\tracking_ms_counter[1]~44_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[1]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[1] .is_wysiwyg = "true";
defparam \tracking_ms_counter[1] .power_up = "low";

dffeas \tracking_ms_counter[4] (
	.clk(clk),
	.d(\tracking_ms_counter[4]~50_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[4]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[4] .is_wysiwyg = "true";
defparam \tracking_ms_counter[4] .power_up = "low";

cycloneiii_lcell_comb \dll_lock_counter[1]~34 (
	.dataa(\dll_lock_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\dll_lock_counter[1]~34_cout ));
defparam \dll_lock_counter[1]~34 .lut_mask = 16'h0055;
defparam \dll_lock_counter[1]~34 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dll_lock_counter[1]~35 (
	.dataa(\dll_lock_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[1]~34_cout ),
	.combout(\dll_lock_counter[1]~35_combout ),
	.cout(\dll_lock_counter[1]~36 ));
defparam \dll_lock_counter[1]~35 .lut_mask = 16'h5AAF;
defparam \dll_lock_counter[1]~35 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[2]~37 (
	.dataa(\dll_lock_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[1]~36 ),
	.combout(\dll_lock_counter[2]~37_combout ),
	.cout(\dll_lock_counter[2]~38 ));
defparam \dll_lock_counter[2]~37 .lut_mask = 16'h5A5F;
defparam \dll_lock_counter[2]~37 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[3]~39 (
	.dataa(\dll_lock_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[2]~38 ),
	.combout(\dll_lock_counter[3]~39_combout ),
	.cout(\dll_lock_counter[3]~40 ));
defparam \dll_lock_counter[3]~39 .lut_mask = 16'h5AAF;
defparam \dll_lock_counter[3]~39 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[4]~41 (
	.dataa(\dll_lock_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[3]~40 ),
	.combout(\dll_lock_counter[4]~41_combout ),
	.cout(\dll_lock_counter[4]~42 ));
defparam \dll_lock_counter[4]~41 .lut_mask = 16'h5A5F;
defparam \dll_lock_counter[4]~41 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[5]~43 (
	.dataa(\dll_lock_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[4]~42 ),
	.combout(\dll_lock_counter[5]~43_combout ),
	.cout(\dll_lock_counter[5]~44 ));
defparam \dll_lock_counter[5]~43 .lut_mask = 16'h5AAF;
defparam \dll_lock_counter[5]~43 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[6]~45 (
	.dataa(\dll_lock_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[5]~44 ),
	.combout(\dll_lock_counter[6]~45_combout ),
	.cout(\dll_lock_counter[6]~46 ));
defparam \dll_lock_counter[6]~45 .lut_mask = 16'h5A5F;
defparam \dll_lock_counter[6]~45 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[7]~47 (
	.dataa(\dll_lock_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[6]~46 ),
	.combout(\dll_lock_counter[7]~47_combout ),
	.cout(\dll_lock_counter[7]~48 ));
defparam \dll_lock_counter[7]~47 .lut_mask = 16'h5AAF;
defparam \dll_lock_counter[7]~47 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[8]~49 (
	.dataa(\dll_lock_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[7]~48 ),
	.combout(\dll_lock_counter[8]~49_combout ),
	.cout(\dll_lock_counter[8]~50 ));
defparam \dll_lock_counter[8]~49 .lut_mask = 16'h5AAF;
defparam \dll_lock_counter[8]~49 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[9]~51 (
	.dataa(\dll_lock_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dll_lock_counter[8]~50 ),
	.combout(\dll_lock_counter[9]~51_combout ),
	.cout(\dll_lock_counter[9]~52 ));
defparam \dll_lock_counter[9]~51 .lut_mask = 16'h5A5F;
defparam \dll_lock_counter[9]~51 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \dll_lock_counter[10]~53 (
	.dataa(\dll_lock_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\dll_lock_counter[9]~52 ),
	.combout(\dll_lock_counter[10]~53_combout ),
	.cout());
defparam \dll_lock_counter[10]~53 .lut_mask = 16'h5A5A;
defparam \dll_lock_counter[10]~53 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \tracking_ms_counter[0]~40 (
	.dataa(\tracking_ms_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\tracking_ms_counter[0]~40_combout ),
	.cout(\tracking_ms_counter[0]~41 ));
defparam \tracking_ms_counter[0]~40 .lut_mask = 16'h55AA;
defparam \tracking_ms_counter[0]~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tracking_ms_counter[1]~44 (
	.dataa(\tracking_ms_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[0]~41 ),
	.combout(\tracking_ms_counter[1]~44_combout ),
	.cout(\tracking_ms_counter[1]~45 ));
defparam \tracking_ms_counter[1]~44 .lut_mask = 16'h5A5F;
defparam \tracking_ms_counter[1]~44 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \tracking_ms_counter[4]~50 (
	.dataa(\tracking_ms_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[3]~49 ),
	.combout(\tracking_ms_counter[4]~50_combout ),
	.cout(\tracking_ms_counter[4]~51 ));
defparam \tracking_ms_counter[4]~50 .lut_mask = 16'h5AAF;
defparam \tracking_ms_counter[4]~50 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~2 (
	.dataa(\milisecond_tick_gen_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~1_cout ),
	.combout(\Add7~2_combout ),
	.cout(\Add7~3 ));
defparam \Add7~2 .lut_mask = 16'h5AAF;
defparam \Add7~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~4 (
	.dataa(\milisecond_tick_gen_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~3 ),
	.combout(\Add7~4_combout ),
	.cout(\Add7~5 ));
defparam \Add7~4 .lut_mask = 16'h5A5F;
defparam \Add7~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~6 (
	.dataa(\milisecond_tick_gen_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~5 ),
	.combout(\Add7~6_combout ),
	.cout(\Add7~7 ));
defparam \Add7~6 .lut_mask = 16'h5A5F;
defparam \Add7~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~8 (
	.dataa(\milisecond_tick_gen_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~7 ),
	.combout(\Add7~8_combout ),
	.cout(\Add7~9 ));
defparam \Add7~8 .lut_mask = 16'h5AAF;
defparam \Add7~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~10 (
	.dataa(\milisecond_tick_gen_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~9 ),
	.combout(\Add7~10_combout ),
	.cout(\Add7~11 ));
defparam \Add7~10 .lut_mask = 16'h5AAF;
defparam \Add7~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~12 (
	.dataa(\milisecond_tick_gen_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~11 ),
	.combout(\Add7~12_combout ),
	.cout(\Add7~13 ));
defparam \Add7~12 .lut_mask = 16'h5A5F;
defparam \Add7~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~14 (
	.dataa(\milisecond_tick_gen_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~13 ),
	.combout(\Add7~14_combout ),
	.cout(\Add7~15 ));
defparam \Add7~14 .lut_mask = 16'h5AAF;
defparam \Add7~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~16 (
	.dataa(\milisecond_tick_gen_count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~15 ),
	.combout(\Add7~16_combout ),
	.cout(\Add7~17 ));
defparam \Add7~16 .lut_mask = 16'h5A5F;
defparam \Add7~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~18 (
	.dataa(\milisecond_tick_gen_count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~17 ),
	.combout(\Add7~18_combout ),
	.cout(\Add7~19 ));
defparam \Add7~18 .lut_mask = 16'h5A5F;
defparam \Add7~18 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~20 (
	.dataa(\milisecond_tick_gen_count[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~19 ),
	.combout(\Add7~20_combout ),
	.cout(\Add7~21 ));
defparam \Add7~20 .lut_mask = 16'h5AAF;
defparam \Add7~20 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~22 (
	.dataa(\milisecond_tick_gen_count[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~21 ),
	.combout(\Add7~22_combout ),
	.cout(\Add7~23 ));
defparam \Add7~22 .lut_mask = 16'h5AAF;
defparam \Add7~22 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~24 (
	.dataa(\milisecond_tick_gen_count[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~23 ),
	.combout(\Add7~24_combout ),
	.cout(\Add7~25 ));
defparam \Add7~24 .lut_mask = 16'h5AAF;
defparam \Add7~24 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~26 (
	.dataa(\milisecond_tick_gen_count[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~25 ),
	.combout(\Add7~26_combout ),
	.cout(\Add7~27 ));
defparam \Add7~26 .lut_mask = 16'h5A5F;
defparam \Add7~26 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~28 (
	.dataa(\milisecond_tick_gen_count[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~27 ),
	.combout(\Add7~28_combout ),
	.cout(\Add7~29 ));
defparam \Add7~28 .lut_mask = 16'h5A5F;
defparam \Add7~28 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~30 (
	.dataa(\milisecond_tick_gen_count[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~29 ),
	.combout(\Add7~30_combout ),
	.cout(\Add7~31 ));
defparam \Add7~30 .lut_mask = 16'h5A5F;
defparam \Add7~30 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~32 (
	.dataa(\milisecond_tick_gen_count[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add7~31 ),
	.combout(\Add7~32_combout ),
	.cout(\Add7~33 ));
defparam \Add7~32 .lut_mask = 16'h5AAF;
defparam \Add7~32 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add7~34 (
	.dataa(\milisecond_tick_gen_count[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add7~33 ),
	.combout(\Add7~34_combout ),
	.cout());
defparam \Add7~34 .lut_mask = 16'h5A5A;
defparam \Add7~34 .sum_lutc_input = "cin";

dffeas \curr_ctrl.command_done (
	.clk(clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_done~q ),
	.prn(vcc));
defparam \curr_ctrl.command_done .is_wysiwyg = "true";
defparam \curr_ctrl.command_done .power_up = "low";

cycloneiii_lcell_comb \Selector1~1 (
	.dataa(admin_ctrlcommand_done),
	.datab(dgwb_ctrlcommand_done),
	.datac(Selector1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector1~2 (
	.dataa(\Selector1~1_combout ),
	.datab(dgrb_ctrlcommand_done),
	.datac(gnd),
	.datad(WideOr11),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hEEFF;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \dll_lock_counter[0] (
	.clk(clk),
	.d(\dll_lock_counter[0]~32_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dll_lock_counter[0]~q ),
	.prn(vcc));
defparam \dll_lock_counter[0] .is_wysiwyg = "true";
defparam \dll_lock_counter[0] .power_up = "low";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\dll_lock_counter[0]~q ),
	.datab(\dll_lock_counter[1]~q ),
	.datac(\dll_lock_counter[2]~q ),
	.datad(\dll_lock_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~1 (
	.dataa(\dll_lock_counter[4]~q ),
	.datab(\dll_lock_counter[5]~q ),
	.datac(\dll_lock_counter[6]~q ),
	.datad(\dll_lock_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFFFE;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~2 (
	.dataa(\dll_lock_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\dll_lock_counter[9]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hAAFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~3 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(\Equal0~2_combout ),
	.datad(\dll_lock_counter[8]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hFF7F;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~0 (
	.dataa(\state.s_operational~q ),
	.datab(\last_state.s_operational~q ),
	.datac(\state.s_prep_customer_mr_setup~q ),
	.datad(curr_cmdcmd_prep_customer_mr_setup),
	.cin(gnd),
	.combout(\WideNor1~0_combout ),
	.cout());
defparam \WideNor1~0 .lut_mask = 16'h6996;
defparam \WideNor1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~1 (
	.dataa(\state.s_write_mtp~q ),
	.datab(curr_cmdcmd_write_mtp),
	.datac(\state.s_was~q ),
	.datad(curr_cmdcmd_was),
	.cin(gnd),
	.combout(\WideNor1~1_combout ),
	.cout());
defparam \WideNor1~1 .lut_mask = 16'h6996;
defparam \WideNor1~1 .sum_lutc_input = "datac";

dffeas \last_state.s_reset (
	.clk(clk),
	.d(\state.s_reset~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_reset~q ),
	.prn(vcc));
defparam \last_state.s_reset .is_wysiwyg = "true";
defparam \last_state.s_reset .power_up = "low";

cycloneiii_lcell_comb \WideNor1~2 (
	.dataa(\state.s_reset~q ),
	.datab(\last_state.s_reset~q ),
	.datac(last_states_rdv),
	.datad(\state.s_rdv~q ),
	.cin(gnd),
	.combout(\WideNor1~2_combout ),
	.cout());
defparam \WideNor1~2 .lut_mask = 16'h6996;
defparam \WideNor1~2 .sum_lutc_input = "datac";

dffeas \last_state.s_cal (
	.clk(clk),
	.d(\state.s_cal~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_cal~q ),
	.prn(vcc));
defparam \last_state.s_cal .is_wysiwyg = "true";
defparam \last_state.s_cal .power_up = "low";

cycloneiii_lcell_comb \WideNor1~3 (
	.dataa(\state.s_cal~q ),
	.datab(\last_state.s_cal~q ),
	.datac(last_states_read_mtp),
	.datad(\state.s_read_mtp~q ),
	.cin(gnd),
	.combout(\WideNor1~3_combout ),
	.cout());
defparam \WideNor1~3 .lut_mask = 16'h6996;
defparam \WideNor1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~4 (
	.dataa(\WideNor1~0_combout ),
	.datab(\WideNor1~1_combout ),
	.datac(\WideNor1~2_combout ),
	.datad(\WideNor1~3_combout ),
	.cin(gnd),
	.combout(\WideNor1~4_combout ),
	.cout());
defparam \WideNor1~4 .lut_mask = 16'hFFFE;
defparam \WideNor1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~5 (
	.dataa(\state.s_phy_initialise~q ),
	.datab(\last_state.s_phy_initialise~q ),
	.datac(\last_state.s_tracking_setup~q ),
	.datad(\state.s_tracking_setup~q ),
	.cin(gnd),
	.combout(\WideNor1~5_combout ),
	.cout());
defparam \WideNor1~5 .lut_mask = 16'h6996;
defparam \WideNor1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal5~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\tracking_ms_counter[0]~q ),
	.datad(\tracking_ms_counter[1]~q ),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'h0FFF;
defparam \Equal5~0 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[17] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[17]~74_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[17]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[17] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[17] .power_up = "low";

dffeas \milisecond_tick_gen_count[14] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[14]~75_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[14]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[14] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[14] .power_up = "low";

dffeas \milisecond_tick_gen_count[16] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[16]~77_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[16]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[16] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[16] .power_up = "low";

dffeas \milisecond_tick_gen_count[15] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[15]~78_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[15]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[15] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[15] .power_up = "low";

cycloneiii_lcell_comb \Equal4~0 (
	.dataa(\milisecond_tick_gen_count[17]~q ),
	.datab(\milisecond_tick_gen_count[14]~q ),
	.datac(\milisecond_tick_gen_count[16]~q ),
	.datad(\milisecond_tick_gen_count[15]~q ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hEFFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[11] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[11]~79_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[11]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[11] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[11] .power_up = "low";

dffeas \milisecond_tick_gen_count[13] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[13]~80_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[13]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[13] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[13] .power_up = "low";

dffeas \milisecond_tick_gen_count[12] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[12]~81_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[12]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[12] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[12] .power_up = "low";

dffeas \milisecond_tick_gen_count[10] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[10]~82_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[10]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[10] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[10] .power_up = "low";

cycloneiii_lcell_comb \Equal4~1 (
	.dataa(\milisecond_tick_gen_count[11]~q ),
	.datab(\milisecond_tick_gen_count[13]~q ),
	.datac(\milisecond_tick_gen_count[12]~q ),
	.datad(\milisecond_tick_gen_count[10]~q ),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
defparam \Equal4~1 .lut_mask = 16'hBFFF;
defparam \Equal4~1 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[8] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[8]~83_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[8]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[8] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[8] .power_up = "low";

dffeas \milisecond_tick_gen_count[7] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[7]~84_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[7]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[7] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[7] .power_up = "low";

dffeas \milisecond_tick_gen_count[6] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[6]~85_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[6]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[6] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[6] .power_up = "low";

dffeas \milisecond_tick_gen_count[9] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[9]~86_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[9]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[9] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[9] .power_up = "low";

cycloneiii_lcell_comb \Equal4~2 (
	.dataa(\milisecond_tick_gen_count[8]~q ),
	.datab(\milisecond_tick_gen_count[7]~q ),
	.datac(\milisecond_tick_gen_count[6]~q ),
	.datad(\milisecond_tick_gen_count[9]~q ),
	.cin(gnd),
	.combout(\Equal4~2_combout ),
	.cout());
defparam \Equal4~2 .lut_mask = 16'hFEFF;
defparam \Equal4~2 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[5] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[5]~87_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[5]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[5] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[5] .power_up = "low";

dffeas \milisecond_tick_gen_count[2] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[2]~88_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[2]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[2] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[2] .power_up = "low";

dffeas \milisecond_tick_gen_count[4] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[4]~89_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[4]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[4] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[4] .power_up = "low";

dffeas \milisecond_tick_gen_count[3] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[3]~90_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[3]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[3] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[3] .power_up = "low";

cycloneiii_lcell_comb \Equal4~3 (
	.dataa(\milisecond_tick_gen_count[5]~q ),
	.datab(\milisecond_tick_gen_count[2]~q ),
	.datac(\milisecond_tick_gen_count[4]~q ),
	.datad(\milisecond_tick_gen_count[3]~q ),
	.cin(gnd),
	.combout(\Equal4~3_combout ),
	.cout());
defparam \Equal4~3 .lut_mask = 16'hEFFF;
defparam \Equal4~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~4 (
	.dataa(\Equal4~0_combout ),
	.datab(\Equal4~1_combout ),
	.datac(\Equal4~2_combout ),
	.datad(\Equal4~3_combout ),
	.cin(gnd),
	.combout(\Equal4~4_combout ),
	.cout());
defparam \Equal4~4 .lut_mask = 16'hFFFE;
defparam \Equal4~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~12 (
	.dataa(\last_state.s_operational~q ),
	.datab(last_states_rdv),
	.datac(\last_state.s_cal~q ),
	.datad(\last_state.s_reset~q ),
	.cin(gnd),
	.combout(\WideNor1~12_combout ),
	.cout());
defparam \WideNor1~12 .lut_mask = 16'hFEFF;
defparam \WideNor1~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dll_lock_counter[0]~32 (
	.dataa(\Equal0~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\dll_lock_counter[0]~q ),
	.cin(gnd),
	.combout(\dll_lock_counter[0]~32_combout ),
	.cout());
defparam \dll_lock_counter[0]~32 .lut_mask = 16'h55FF;
defparam \dll_lock_counter[0]~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[17]~74 (
	.dataa(\milisecond_tick_gen_count[17]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~34_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[17]~74_combout ),
	.cout());
defparam \milisecond_tick_gen_count[17]~74 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[17]~74 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[14]~75 (
	.dataa(\milisecond_tick_gen_count[14]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~28_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[14]~75_combout ),
	.cout());
defparam \milisecond_tick_gen_count[14]~75 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[14]~75 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[0]~76 (
	.dataa(\state.s_operational~q ),
	.datab(\last_state.s_operational~q ),
	.datac(gnd),
	.datad(\Equal4~5_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[0]~76_combout ),
	.cout());
defparam \milisecond_tick_gen_count[0]~76 .lut_mask = 16'hEEFF;
defparam \milisecond_tick_gen_count[0]~76 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[16]~77 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~32_combout ),
	.datac(\milisecond_tick_gen_count[16]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[16]~77_combout ),
	.cout());
defparam \milisecond_tick_gen_count[16]~77 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[16]~77 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[15]~78 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~30_combout ),
	.datac(\milisecond_tick_gen_count[15]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[15]~78_combout ),
	.cout());
defparam \milisecond_tick_gen_count[15]~78 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[15]~78 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[11]~79 (
	.dataa(\milisecond_tick_gen_count[11]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~22_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[11]~79_combout ),
	.cout());
defparam \milisecond_tick_gen_count[11]~79 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[11]~79 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[13]~80 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~26_combout ),
	.datac(\milisecond_tick_gen_count[13]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[13]~80_combout ),
	.cout());
defparam \milisecond_tick_gen_count[13]~80 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[13]~80 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[12]~81 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~24_combout ),
	.datac(\milisecond_tick_gen_count[12]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[12]~81_combout ),
	.cout());
defparam \milisecond_tick_gen_count[12]~81 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[12]~81 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[10]~82 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~20_combout ),
	.datac(\milisecond_tick_gen_count[10]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[10]~82_combout ),
	.cout());
defparam \milisecond_tick_gen_count[10]~82 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[10]~82 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[8]~83 (
	.dataa(\milisecond_tick_gen_count[8]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~16_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[8]~83_combout ),
	.cout());
defparam \milisecond_tick_gen_count[8]~83 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[8]~83 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[7]~84 (
	.dataa(\milisecond_tick_gen_count[7]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~14_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[7]~84_combout ),
	.cout());
defparam \milisecond_tick_gen_count[7]~84 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[7]~84 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[6]~85 (
	.dataa(\milisecond_tick_gen_count[6]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~12_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[6]~85_combout ),
	.cout());
defparam \milisecond_tick_gen_count[6]~85 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[6]~85 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[9]~86 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~18_combout ),
	.datac(\milisecond_tick_gen_count[9]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[9]~86_combout ),
	.cout());
defparam \milisecond_tick_gen_count[9]~86 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[9]~86 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[5]~87 (
	.dataa(\milisecond_tick_gen_count[5]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~10_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[5]~87_combout ),
	.cout());
defparam \milisecond_tick_gen_count[5]~87 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[5]~87 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[2]~88 (
	.dataa(\milisecond_tick_gen_count[2]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~4_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[2]~88_combout ),
	.cout());
defparam \milisecond_tick_gen_count[2]~88 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[2]~88 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[4]~89 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~8_combout ),
	.datac(\milisecond_tick_gen_count[4]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[4]~89_combout ),
	.cout());
defparam \milisecond_tick_gen_count[4]~89 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[4]~89 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[3]~90 (
	.dataa(\milisecond_tick_gen_count[0]~76_combout ),
	.datab(\Add7~6_combout ),
	.datac(\milisecond_tick_gen_count[3]~q ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[3]~90_combout ),
	.cout());
defparam \milisecond_tick_gen_count[3]~90 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[3]~90 .sum_lutc_input = "datac";

dffeas \mtp_almt:dvw_size_a0[5] (
	.clk(clk),
	.d(\curr_ctrl.command_result[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[5]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[5] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[5] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[4] (
	.clk(clk),
	.d(\curr_ctrl.command_result[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[4]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[4] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[4] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[3] (
	.clk(clk),
	.d(\curr_ctrl.command_result[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[3]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[3] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[3] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[2] (
	.clk(clk),
	.d(\curr_ctrl.command_result[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[2]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[2] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[2] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[1] (
	.clk(clk),
	.d(\curr_ctrl.command_result[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[1]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[1] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[1] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[0] (
	.clk(clk),
	.d(\curr_ctrl.command_result[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a0[0]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[0] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[0] .power_up = "low";

cycloneiii_lcell_comb \mtp_almt:dvw_size_a0[0]~0 (
	.dataa(\curr_ctrl.command_done~q ),
	.datab(\state.s_read_mtp~q ),
	.datac(\mtp_almts_checked[1]~q ),
	.datad(\mtp_almts_checked[0]~q ),
	.cin(gnd),
	.combout(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.cout());
defparam \mtp_almt:dvw_size_a0[0]~0 .lut_mask = 16'hEFFF;
defparam \mtp_almt:dvw_size_a0[0]~0 .sum_lutc_input = "datac";

dffeas ctl_init_success(
	.clk(clk),
	.d(\int_ctl_init_success~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_success1),
	.prn(vcc));
defparam ctl_init_success.is_wysiwyg = "true";
defparam ctl_init_success.power_up = "low";

dffeas \state.s_init_dram (
	.clk(clk),
	.d(\state.s_phy_initialise~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(states_init_dram),
	.prn(vcc));
defparam \state.s_init_dram .is_wysiwyg = "true";
defparam \state.s_init_dram .power_up = "low";

cycloneiii_lcell_comb \WideOr34~8 (
	.dataa(\WideOr34~6_combout ),
	.datab(\WideOr34~7_combout ),
	.datac(gnd),
	.datad(\state.s_prep_customer_mr_setup~q ),
	.cin(gnd),
	.combout(WideOr34),
	.cout());
defparam \WideOr34~8 .lut_mask = 16'hEEFF;
defparam \WideOr34~8 .sum_lutc_input = "datac";

dffeas \curr_cmd.cmd_prep_customer_mr_setup (
	.clk(clk),
	.d(\state.s_prep_customer_mr_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_prep_customer_mr_setup),
	.prn(vcc));
defparam \curr_cmd.cmd_prep_customer_mr_setup .is_wysiwyg = "true";
defparam \curr_cmd.cmd_prep_customer_mr_setup .power_up = "low";

cycloneiii_lcell_comb \Selector1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datad(curr_cmdcmd_prep_customer_mr_setup),
	.cin(gnd),
	.combout(Selector1),
	.cout());
defparam \Selector1~0 .lut_mask = 16'h0FFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \curr_cmd.cmd_write_btp (
	.clk(clk),
	.d(\state.s_write_btp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_write_btp),
	.prn(vcc));
defparam \curr_cmd.cmd_write_btp .is_wysiwyg = "true";
defparam \curr_cmd.cmd_write_btp .power_up = "low";

dffeas \curr_cmd.cmd_write_mtp (
	.clk(clk),
	.d(\state.s_write_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_write_mtp),
	.prn(vcc));
defparam \curr_cmd.cmd_write_mtp .is_wysiwyg = "true";
defparam \curr_cmd.cmd_write_mtp .power_up = "low";

dffeas \curr_cmd.cmd_was (
	.clk(clk),
	.d(\state.s_was~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_was),
	.prn(vcc));
defparam \curr_cmd.cmd_was .is_wysiwyg = "true";
defparam \curr_cmd.cmd_was .power_up = "low";

cycloneiii_lcell_comb \WideOr0~0 (
	.dataa(gnd),
	.datab(curr_cmdcmd_write_btp),
	.datac(curr_cmdcmd_write_mtp),
	.datad(curr_cmdcmd_was),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'h3FFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

dffeas \curr_cmd.cmd_idle (
	.clk(clk),
	.d(\Selector41~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_idle),
	.prn(vcc));
defparam \curr_cmd.cmd_idle .is_wysiwyg = "true";
defparam \curr_cmd.cmd_idle .power_up = "low";

cycloneiii_lcell_comb WideOr1(
	.dataa(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datab(curr_cmdcmd_prep_customer_mr_setup),
	.datac(curr_cmdcmd_idle),
	.datad(WideOr0),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hEFFF;
defparam WideOr1.sum_lutc_input = "datac";

dffeas \last_state.s_rdv (
	.clk(clk),
	.d(\state.s_rdv~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_rdv),
	.prn(vcc));
defparam \last_state.s_rdv .is_wysiwyg = "true";
defparam \last_state.s_rdv .power_up = "low";

dffeas \last_state.s_read_mtp (
	.clk(clk),
	.d(\state.s_read_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_read_mtp),
	.prn(vcc));
defparam \last_state.s_read_mtp .is_wysiwyg = "true";
defparam \last_state.s_read_mtp .power_up = "low";

dffeas \last_state.s_rrp_seek (
	.clk(clk),
	.d(\state.s_rrp_seek~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_rrp_seek),
	.prn(vcc));
defparam \last_state.s_rrp_seek .is_wysiwyg = "true";
defparam \last_state.s_rrp_seek .power_up = "low";

dffeas \last_state.s_adv_rd_lat (
	.clk(clk),
	.d(\state.s_adv_rd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_adv_rd_lat),
	.prn(vcc));
defparam \last_state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \last_state.s_adv_rd_lat .power_up = "low";

dffeas \last_state.s_rrp_sweep (
	.clk(clk),
	.d(\state.s_rrp_sweep~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_rrp_sweep),
	.prn(vcc));
defparam \last_state.s_rrp_sweep .is_wysiwyg = "true";
defparam \last_state.s_rrp_sweep .power_up = "low";

dffeas \last_state.s_adv_wr_lat (
	.clk(clk),
	.d(\state.s_adv_wr_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_adv_wr_lat),
	.prn(vcc));
defparam \last_state.s_adv_wr_lat .is_wysiwyg = "true";
defparam \last_state.s_adv_wr_lat .power_up = "low";

dffeas \last_state.s_rrp_reset (
	.clk(clk),
	.d(\state.s_rrp_reset~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(last_states_rrp_reset),
	.prn(vcc));
defparam \last_state.s_rrp_reset .is_wysiwyg = "true";
defparam \last_state.s_rrp_reset .power_up = "low";

cycloneiii_lcell_comb \Selector58~0 (
	.dataa(\WideOr34~6_combout ),
	.datab(\WideNor1~11_combout ),
	.datac(gnd),
	.datad(\state.s_poa~q ),
	.cin(gnd),
	.combout(Selector58),
	.cout());
defparam \Selector58~0 .lut_mask = 16'hEEFF;
defparam \Selector58~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ctrl_op_rec.command_op.single_bit~0 (
	.dataa(\state.s_read_mtp~q ),
	.datab(\state.s_rrp_sweep~q ),
	.datac(\state.s_poa~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(ctrl_op_reccommand_opsingle_bit),
	.cout());
defparam \ctrl_op_rec.command_op.single_bit~0 .lut_mask = 16'hFEFE;
defparam \ctrl_op_rec.command_op.single_bit~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ctrl_op_rec.command_op.mtp_almt~0 (
	.dataa(ctrl_op_reccommand_opsingle_bit),
	.datab(\mtp_almts_checked[0]~q ),
	.datac(\mtp_almts_checked[1]~q ),
	.datad(\mtp_correct_almt~q ),
	.cin(gnd),
	.combout(ctrl_op_reccommand_opmtp_almt),
	.cout());
defparam \ctrl_op_rec.command_op.mtp_almt~0 .lut_mask = 16'hFFFE;
defparam \ctrl_op_rec.command_op.mtp_almt~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector57~0 (
	.dataa(\WideOr34~6_combout ),
	.datab(\master_ctrl_op_rec~41_combout ),
	.datac(\state.s_tracking~q ),
	.datad(\state.s_tracking_setup~q ),
	.cin(gnd),
	.combout(Selector57),
	.cout());
defparam \Selector57~0 .lut_mask = 16'hFFFE;
defparam \Selector57~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector52~0 (
	.dataa(\state.s_poa~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\WideNor1~16_combout ),
	.cin(gnd),
	.combout(Selector52),
	.cout());
defparam \Selector52~0 .lut_mask = 16'hAAFF;
defparam \Selector52~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tracking_ms_counter[2]~46 (
	.dataa(\tracking_ms_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[1]~45 ),
	.combout(\tracking_ms_counter[2]~46_combout ),
	.cout(\tracking_ms_counter[2]~47 ));
defparam \tracking_ms_counter[2]~46 .lut_mask = 16'h5AAF;
defparam \tracking_ms_counter[2]~46 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \tracking_ms_counter[3]~48 (
	.dataa(\tracking_ms_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[2]~47 ),
	.combout(\tracking_ms_counter[3]~48_combout ),
	.cout(\tracking_ms_counter[3]~49 ));
defparam \tracking_ms_counter[3]~48 .lut_mask = 16'h5A5F;
defparam \tracking_ms_counter[3]~48 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \tracking_ms_counter[5]~52 (
	.dataa(\tracking_ms_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[4]~51 ),
	.combout(\tracking_ms_counter[5]~52_combout ),
	.cout(\tracking_ms_counter[5]~53 ));
defparam \tracking_ms_counter[5]~52 .lut_mask = 16'h5A5F;
defparam \tracking_ms_counter[5]~52 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Selector34~0 (
	.dataa(\state.s_read_mtp~q ),
	.datab(gnd),
	.datac(\mtp_almts_checked[1]~q ),
	.datad(\mtp_almts_checked[0]~q ),
	.cin(gnd),
	.combout(\Selector34~0_combout ),
	.cout());
defparam \Selector34~0 .lut_mask = 16'hAFFF;
defparam \Selector34~0 .sum_lutc_input = "datac";

dffeas \last_state.s_tracking (
	.clk(clk),
	.d(\state.s_tracking~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_tracking~q ),
	.prn(vcc));
defparam \last_state.s_tracking .is_wysiwyg = "true";
defparam \last_state.s_tracking .power_up = "low";

cycloneiii_lcell_comb \WideNor1~6 (
	.dataa(\state.s_tracking~q ),
	.datab(\last_state.s_tracking~q ),
	.datac(last_states_rrp_seek),
	.datad(\state.s_rrp_seek~q ),
	.cin(gnd),
	.combout(\WideNor1~6_combout ),
	.cout());
defparam \WideNor1~6 .lut_mask = 16'h6996;
defparam \WideNor1~6 .sum_lutc_input = "datac";

dffeas \state.s_write_btp (
	.clk(clk),
	.d(\state.s_cal~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_write_btp~q ),
	.prn(vcc));
defparam \state.s_write_btp .is_wysiwyg = "true";
defparam \state.s_write_btp .power_up = "low";

cycloneiii_lcell_comb \WideNor1~7 (
	.dataa(states_init_dram),
	.datab(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datac(\state.s_write_btp~q ),
	.datad(curr_cmdcmd_write_btp),
	.cin(gnd),
	.combout(\WideNor1~7_combout ),
	.cout());
defparam \WideNor1~7 .lut_mask = 16'h6996;
defparam \WideNor1~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state~163 (
	.dataa(\mtp_almts_checked[1]~q ),
	.datab(gnd),
	.datac(\mtp_almts_checked[0]~q ),
	.datad(\state.s_rrp_sweep~q ),
	.cin(gnd),
	.combout(\state~163_combout ),
	.cout());
defparam \state~163 .lut_mask = 16'hFFF5;
defparam \state~163 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \hold_state~2 (
	.dataa(\state~162_combout ),
	.datab(\tracking_update_due~q ),
	.datac(gnd),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\hold_state~2_combout ),
	.cout());
defparam \hold_state~2 .lut_mask = 16'hEEFF;
defparam \hold_state~2 .sum_lutc_input = "datac";

dffeas \state.s_read_mtp (
	.clk(clk),
	.d(\state~163_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\hold_state~2_combout ),
	.q(\state.s_read_mtp~q ),
	.prn(vcc));
defparam \state.s_read_mtp .is_wysiwyg = "true";
defparam \state.s_read_mtp .power_up = "low";

cycloneiii_lcell_comb \state~46 (
	.dataa(\state.s_write_mtp~q ),
	.datab(\state.s_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~46_combout ),
	.cout());
defparam \state~46 .lut_mask = 16'hEEEE;
defparam \state~46 .sum_lutc_input = "datac";

dffeas \state.s_rrp_reset (
	.clk(clk),
	.d(\state~46_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_rrp_reset~q ),
	.prn(vcc));
defparam \state.s_rrp_reset .is_wysiwyg = "true";
defparam \state.s_rrp_reset .power_up = "low";

dffeas \state.s_rrp_sweep (
	.clk(clk),
	.d(\state.s_rrp_reset~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_rrp_sweep~q ),
	.prn(vcc));
defparam \state.s_rrp_sweep .is_wysiwyg = "true";
defparam \state.s_rrp_sweep .power_up = "low";

cycloneiii_lcell_comb \WideNor1~8 (
	.dataa(last_states_adv_rd_lat),
	.datab(\state.s_adv_rd_lat~q ),
	.datac(last_states_rrp_sweep),
	.datad(\state.s_rrp_sweep~q ),
	.cin(gnd),
	.combout(\WideNor1~8_combout ),
	.cout());
defparam \WideNor1~8 .lut_mask = 16'h6996;
defparam \WideNor1~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~9 (
	.dataa(\WideNor1~5_combout ),
	.datab(\WideNor1~6_combout ),
	.datac(\WideNor1~7_combout ),
	.datad(\WideNor1~8_combout ),
	.cin(gnd),
	.combout(\WideNor1~9_combout ),
	.cout());
defparam \WideNor1~9 .lut_mask = 16'hFFFE;
defparam \WideNor1~9 .sum_lutc_input = "datac";

dffeas \last_state.s_poa (
	.clk(clk),
	.d(\state.s_poa~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_poa~q ),
	.prn(vcc));
defparam \last_state.s_poa .is_wysiwyg = "true";
defparam \last_state.s_poa .power_up = "low";

cycloneiii_lcell_comb \WideNor1~10 (
	.dataa(\state.s_poa~q ),
	.datab(\last_state.s_poa~q ),
	.datac(last_states_adv_wr_lat),
	.datad(\state.s_adv_wr_lat~q ),
	.cin(gnd),
	.combout(\WideNor1~10_combout ),
	.cout());
defparam \WideNor1~10 .lut_mask = 16'h6996;
defparam \WideNor1~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \process_14~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(last_states_rrp_reset),
	.datad(\state.s_rrp_reset~q ),
	.cin(gnd),
	.combout(\process_14~13_combout ),
	.cout());
defparam \process_14~13 .lut_mask = 16'h0FF0;
defparam \process_14~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~11 (
	.dataa(\WideNor1~4_combout ),
	.datab(\WideNor1~9_combout ),
	.datac(\WideNor1~10_combout ),
	.datad(\process_14~13_combout ),
	.cin(gnd),
	.combout(\WideNor1~11_combout ),
	.cout());
defparam \WideNor1~11 .lut_mask = 16'hFFFE;
defparam \WideNor1~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr28~0 (
	.dataa(\state.s_reset~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\WideOr28~0_combout ),
	.cout());
defparam \WideOr28~0 .lut_mask = 16'hAAFF;
defparam \WideOr28~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dis_state~5 (
	.dataa(\state.s_cal~q ),
	.datab(\dis_state~q ),
	.datac(\WideNor1~11_combout ),
	.datad(\WideOr28~0_combout ),
	.cin(gnd),
	.combout(\dis_state~5_combout ),
	.cout());
defparam \dis_state~5 .lut_mask = 16'hEFFF;
defparam \dis_state~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \master_ctrl_op_rec~41 (
	.dataa(\state.s_reset~q ),
	.datab(\state.s_operational~q ),
	.datac(\state.s_poa~q ),
	.datad(\WideNor1~11_combout ),
	.cin(gnd),
	.combout(\master_ctrl_op_rec~41_combout ),
	.cout());
defparam \master_ctrl_op_rec~41 .lut_mask = 16'hBFFF;
defparam \master_ctrl_op_rec~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \state.s_phy_initialise~1 (
	.dataa(\state.s_reset~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state.s_phy_initialise~1_combout ),
	.cout());
defparam \state.s_phy_initialise~1 .lut_mask = 16'h5555;
defparam \state.s_phy_initialise~1 .sum_lutc_input = "datac";

dffeas \state.s_phy_initialise (
	.clk(clk),
	.d(\state.s_phy_initialise~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_phy_initialise~q ),
	.prn(vcc));
defparam \state.s_phy_initialise .is_wysiwyg = "true";
defparam \state.s_phy_initialise .power_up = "low";

cycloneiii_lcell_comb \dis_state~6 (
	.dataa(\Equal0~3_combout ),
	.datab(\dis_state~5_combout ),
	.datac(\master_ctrl_op_rec~41_combout ),
	.datad(\state.s_phy_initialise~q ),
	.cin(gnd),
	.combout(\dis_state~6_combout ),
	.cout());
defparam \dis_state~6 .lut_mask = 16'hCF5F;
defparam \dis_state~6 .sum_lutc_input = "datac";

dffeas dis_state(
	.clk(clk),
	.d(\dis_state~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dis_state~q ),
	.prn(vcc));
defparam dis_state.is_wysiwyg = "true";
defparam dis_state.power_up = "low";

dffeas hold_state(
	.clk(clk),
	.d(\hold_state~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hold_state~q ),
	.prn(vcc));
defparam hold_state.is_wysiwyg = "true";
defparam hold_state.power_up = "low";

cycloneiii_lcell_comb \state~162 (
	.dataa(\curr_ctrl.command_done~q ),
	.datab(\dis_state~q ),
	.datac(gnd),
	.datad(\hold_state~q ),
	.cin(gnd),
	.combout(\state~162_combout ),
	.cout());
defparam \state~162 .lut_mask = 16'hEEFF;
defparam \state~162 .sum_lutc_input = "datac";

dffeas \state.s_cal (
	.clk(clk),
	.d(states_init_dram),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_cal~q ),
	.prn(vcc));
defparam \state.s_cal .is_wysiwyg = "true";
defparam \state.s_cal .power_up = "low";

cycloneiii_lcell_comb \mtp_almts_checked[1]~8 (
	.dataa(\state~162_combout ),
	.datab(\state.s_cal~q ),
	.datac(\state.s_read_mtp~q ),
	.datad(\state.s_adv_wr_lat~q ),
	.cin(gnd),
	.combout(\mtp_almts_checked[1]~8_combout ),
	.cout());
defparam \mtp_almts_checked[1]~8 .lut_mask = 16'hFEFF;
defparam \mtp_almts_checked[1]~8 .sum_lutc_input = "datac";

dffeas \mtp_almts_checked[0] (
	.clk(clk),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almts_checked[1]~8_combout ),
	.q(\mtp_almts_checked[0]~q ),
	.prn(vcc));
defparam \mtp_almts_checked[0] .is_wysiwyg = "true";
defparam \mtp_almts_checked[0] .power_up = "low";

cycloneiii_lcell_comb \Selector33~0 (
	.dataa(\state.s_read_mtp~q ),
	.datab(gnd),
	.datac(\mtp_almts_checked[1]~q ),
	.datad(\mtp_almts_checked[0]~q ),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'hAFFA;
defparam \Selector33~0 .sum_lutc_input = "datac";

dffeas \mtp_almts_checked[1] (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almts_checked[1]~8_combout ),
	.q(\mtp_almts_checked[1]~q ),
	.prn(vcc));
defparam \mtp_almts_checked[1] .is_wysiwyg = "true";
defparam \mtp_almts_checked[1] .power_up = "low";

cycloneiii_lcell_comb \state~164 (
	.dataa(\state.s_rrp_sweep~q ),
	.datab(\mtp_almts_checked[1]~q ),
	.datac(gnd),
	.datad(\mtp_almts_checked[0]~q ),
	.cin(gnd),
	.combout(\state~164_combout ),
	.cout());
defparam \state~164 .lut_mask = 16'hEEFF;
defparam \state~164 .sum_lutc_input = "datac";

dffeas \state.s_rrp_seek (
	.clk(clk),
	.d(\state~164_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\hold_state~2_combout ),
	.q(\state.s_rrp_seek~q ),
	.prn(vcc));
defparam \state.s_rrp_seek .is_wysiwyg = "true";
defparam \state.s_rrp_seek .power_up = "low";

dffeas \state.s_rdv (
	.clk(clk),
	.d(\state.s_rrp_seek~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_rdv~q ),
	.prn(vcc));
defparam \state.s_rdv .is_wysiwyg = "true";
defparam \state.s_rdv .power_up = "low";

dffeas \state.s_was (
	.clk(clk),
	.d(\state.s_rdv~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_was~q ),
	.prn(vcc));
defparam \state.s_was .is_wysiwyg = "true";
defparam \state.s_was .power_up = "low";

dffeas \state.s_adv_rd_lat (
	.clk(clk),
	.d(\state.s_was~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_adv_rd_lat~q ),
	.prn(vcc));
defparam \state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \state.s_adv_rd_lat .power_up = "low";

dffeas \state.s_adv_wr_lat (
	.clk(clk),
	.d(\state.s_adv_rd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_adv_wr_lat~q ),
	.prn(vcc));
defparam \state.s_adv_wr_lat .is_wysiwyg = "true";
defparam \state.s_adv_wr_lat .power_up = "low";

dffeas \state.s_poa (
	.clk(clk),
	.d(\state.s_adv_wr_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_poa~q ),
	.prn(vcc));
defparam \state.s_poa .is_wysiwyg = "true";
defparam \state.s_poa .power_up = "low";

dffeas \state.s_tracking_setup (
	.clk(clk),
	.d(\state.s_poa~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_tracking_setup~q ),
	.prn(vcc));
defparam \state.s_tracking_setup .is_wysiwyg = "true";
defparam \state.s_tracking_setup .power_up = "low";

dffeas \state.s_prep_customer_mr_setup (
	.clk(clk),
	.d(\state.s_tracking_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_prep_customer_mr_setup~q ),
	.prn(vcc));
defparam \state.s_prep_customer_mr_setup .is_wysiwyg = "true";
defparam \state.s_prep_customer_mr_setup .power_up = "low";

cycloneiii_lcell_comb \Selector30~0 (
	.dataa(\state.s_tracking~q ),
	.datab(\state.s_prep_customer_mr_setup~q ),
	.datac(\state.s_operational~q ),
	.datad(\tracking_update_due~q ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
defparam \Selector30~0 .lut_mask = 16'hFEFF;
defparam \Selector30~0 .sum_lutc_input = "datac";

dffeas \state.s_operational (
	.clk(clk),
	.d(\Selector30~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_operational~q ),
	.prn(vcc));
defparam \state.s_operational .is_wysiwyg = "true";
defparam \state.s_operational .power_up = "low";

dffeas \last_state.s_operational (
	.clk(clk),
	.d(\state.s_operational~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_operational~q ),
	.prn(vcc));
defparam \last_state.s_operational .is_wysiwyg = "true";
defparam \last_state.s_operational .power_up = "low";

cycloneiii_lcell_comb \process_16~0 (
	.dataa(\state.s_operational~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\last_state.s_operational~q ),
	.cin(gnd),
	.combout(\process_16~0_combout ),
	.cout());
defparam \process_16~0 .lut_mask = 16'hAAFF;
defparam \process_16~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[0]~73 (
	.dataa(\tracking_update_due~q ),
	.datab(\last_state.s_operational~q ),
	.datac(\state.s_operational~q ),
	.datad(\Equal4~5_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[0]~73_combout ),
	.cout());
defparam \milisecond_tick_gen_count[0]~73 .lut_mask = 16'hEFFF;
defparam \milisecond_tick_gen_count[0]~73 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[0]~92 (
	.dataa(\milisecond_tick_gen_count[0]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[0]~92_combout ),
	.cout());
defparam \milisecond_tick_gen_count[0]~92 .lut_mask = 16'hF6F6;
defparam \milisecond_tick_gen_count[0]~92 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[0] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[0]~92_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[0]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[0] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[0] .power_up = "low";

cycloneiii_lcell_comb \Equal4~5 (
	.dataa(\Equal4~4_combout ),
	.datab(\milisecond_tick_gen_count[1]~q ),
	.datac(\milisecond_tick_gen_count[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal4~5_combout ),
	.cout());
defparam \Equal4~5 .lut_mask = 16'hFEFE;
defparam \Equal4~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[2]~72 (
	.dataa(\tracking_update_due~q ),
	.datab(\last_state.s_operational~q ),
	.datac(\Equal4~5_combout ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[2]~72_combout ),
	.cout());
defparam \milisecond_tick_gen_count[2]~72 .lut_mask = 16'hFEFF;
defparam \milisecond_tick_gen_count[2]~72 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add7~1 (
	.dataa(\milisecond_tick_gen_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add7~1_cout ));
defparam \Add7~1 .lut_mask = 16'h0055;
defparam \Add7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \milisecond_tick_gen_count[1]~91 (
	.dataa(\milisecond_tick_gen_count[1]~q ),
	.datab(\milisecond_tick_gen_count[2]~72_combout ),
	.datac(\milisecond_tick_gen_count[0]~73_combout ),
	.datad(\Add7~2_combout ),
	.cin(gnd),
	.combout(\milisecond_tick_gen_count[1]~91_combout ),
	.cout());
defparam \milisecond_tick_gen_count[1]~91 .lut_mask = 16'hB8FF;
defparam \milisecond_tick_gen_count[1]~91 .sum_lutc_input = "datac";

dffeas \milisecond_tick_gen_count[1] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[1]~91_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\milisecond_tick_gen_count[1]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[1] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[1] .power_up = "low";

cycloneiii_lcell_comb \tracking_ms_counter[0]~42 (
	.dataa(\Equal4~4_combout ),
	.datab(\milisecond_tick_gen_count[1]~q ),
	.datac(\milisecond_tick_gen_count[0]~q ),
	.datad(\tracking_update_due~q ),
	.cin(gnd),
	.combout(\tracking_ms_counter[0]~42_combout ),
	.cout());
defparam \tracking_ms_counter[0]~42 .lut_mask = 16'hFEFF;
defparam \tracking_ms_counter[0]~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tracking_ms_counter[0]~43 (
	.dataa(\last_state.s_operational~q ),
	.datab(\Equal5~2_combout ),
	.datac(\tracking_ms_counter[0]~42_combout ),
	.datad(\state.s_operational~q ),
	.cin(gnd),
	.combout(\tracking_ms_counter[0]~43_combout ),
	.cout());
defparam \tracking_ms_counter[0]~43 .lut_mask = 16'hFFF7;
defparam \tracking_ms_counter[0]~43 .sum_lutc_input = "datac";

dffeas \tracking_ms_counter[5] (
	.clk(clk),
	.d(\tracking_ms_counter[5]~52_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[5]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[5] .is_wysiwyg = "true";
defparam \tracking_ms_counter[5] .power_up = "low";

cycloneiii_lcell_comb \tracking_ms_counter[6]~54 (
	.dataa(\tracking_ms_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tracking_ms_counter[5]~53 ),
	.combout(\tracking_ms_counter[6]~54_combout ),
	.cout(\tracking_ms_counter[6]~55 ));
defparam \tracking_ms_counter[6]~54 .lut_mask = 16'h5AAF;
defparam \tracking_ms_counter[6]~54 .sum_lutc_input = "cin";

dffeas \tracking_ms_counter[6] (
	.clk(clk),
	.d(\tracking_ms_counter[6]~54_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[6]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[6] .is_wysiwyg = "true";
defparam \tracking_ms_counter[6] .power_up = "low";

cycloneiii_lcell_comb \tracking_ms_counter[7]~56 (
	.dataa(\tracking_ms_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\tracking_ms_counter[6]~55 ),
	.combout(\tracking_ms_counter[7]~56_combout ),
	.cout());
defparam \tracking_ms_counter[7]~56 .lut_mask = 16'h5A5A;
defparam \tracking_ms_counter[7]~56 .sum_lutc_input = "cin";

dffeas \tracking_ms_counter[7] (
	.clk(clk),
	.d(\tracking_ms_counter[7]~56_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[7]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[7] .is_wysiwyg = "true";
defparam \tracking_ms_counter[7] .power_up = "low";

cycloneiii_lcell_comb \Equal5~1 (
	.dataa(\tracking_ms_counter[4]~q ),
	.datab(\tracking_ms_counter[5]~q ),
	.datac(\tracking_ms_counter[6]~q ),
	.datad(\tracking_ms_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'h7FFF;
defparam \Equal5~1 .sum_lutc_input = "datac";

dffeas \tracking_ms_counter[2] (
	.clk(clk),
	.d(\tracking_ms_counter[2]~46_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[2]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[2] .is_wysiwyg = "true";
defparam \tracking_ms_counter[2] .power_up = "low";

dffeas \tracking_ms_counter[3] (
	.clk(clk),
	.d(\tracking_ms_counter[3]~48_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~43_combout ),
	.q(\tracking_ms_counter[3]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[3] .is_wysiwyg = "true";
defparam \tracking_ms_counter[3] .power_up = "low";

cycloneiii_lcell_comb \Equal5~2 (
	.dataa(\Equal5~0_combout ),
	.datab(\Equal5~1_combout ),
	.datac(\tracking_ms_counter[2]~q ),
	.datad(\tracking_ms_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal5~2_combout ),
	.cout());
defparam \Equal5~2 .lut_mask = 16'hEFFF;
defparam \Equal5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \tracking_update_due~5 (
	.dataa(\tracking_update_due~q ),
	.datab(\Equal5~2_combout ),
	.datac(\Equal4~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\tracking_update_due~5_combout ),
	.cout());
defparam \tracking_update_due~5 .lut_mask = 16'hFEFE;
defparam \tracking_update_due~5 .sum_lutc_input = "datac";

dffeas tracking_update_due(
	.clk(clk),
	.d(\tracking_update_due~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\state.s_operational~q ),
	.sload(gnd),
	.ena(!\process_16~0_combout ),
	.q(\tracking_update_due~q ),
	.prn(vcc));
defparam tracking_update_due.is_wysiwyg = "true";
defparam tracking_update_due.power_up = "low";

cycloneiii_lcell_comb \Selector29~0 (
	.dataa(\state.s_operational~q ),
	.datab(\tracking_update_due~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
defparam \Selector29~0 .lut_mask = 16'hEEEE;
defparam \Selector29~0 .sum_lutc_input = "datac";

dffeas \state.s_tracking (
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_tracking~q ),
	.prn(vcc));
defparam \state.s_tracking .is_wysiwyg = "true";
defparam \state.s_tracking .power_up = "low";

cycloneiii_lcell_comb \Selector37~0 (
	.dataa(\state.s_operational~q ),
	.datab(\int_ctl_init_success~q ),
	.datac(\state.s_tracking~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector37~0_combout ),
	.cout());
defparam \Selector37~0 .lut_mask = 16'hFEFE;
defparam \Selector37~0 .sum_lutc_input = "datac";

dffeas int_ctl_init_success(
	.clk(clk),
	.d(\Selector37~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\int_ctl_init_success~q ),
	.prn(vcc));
defparam int_ctl_init_success.is_wysiwyg = "true";
defparam int_ctl_init_success.power_up = "low";

dffeas \state.s_reset (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_reset~q ),
	.prn(vcc));
defparam \state.s_reset .is_wysiwyg = "true";
defparam \state.s_reset .power_up = "low";

cycloneiii_lcell_comb \WideOr34~6 (
	.dataa(\state.s_reset~q ),
	.datab(\state.s_operational~q ),
	.datac(\state.s_phy_initialise~q ),
	.datad(\state.s_cal~q ),
	.cin(gnd),
	.combout(\WideOr34~6_combout ),
	.cout());
defparam \WideOr34~6 .lut_mask = 16'hBFFF;
defparam \WideOr34~6 .sum_lutc_input = "datac";

dffeas \state.s_write_mtp (
	.clk(clk),
	.d(\state.s_write_btp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~162_combout ),
	.q(\state.s_write_mtp~q ),
	.prn(vcc));
defparam \state.s_write_mtp .is_wysiwyg = "true";
defparam \state.s_write_mtp .power_up = "low";

cycloneiii_lcell_comb \WideOr34~7 (
	.dataa(states_init_dram),
	.datab(\state.s_write_btp~q ),
	.datac(\state.s_write_mtp~q ),
	.datad(\state.s_was~q ),
	.cin(gnd),
	.combout(\WideOr34~7_combout ),
	.cout());
defparam \WideOr34~7 .lut_mask = 16'h7FFF;
defparam \WideOr34~7 .sum_lutc_input = "datac";

dffeas \last_state.s_tracking_setup (
	.clk(clk),
	.d(\state.s_tracking_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_tracking_setup~q ),
	.prn(vcc));
defparam \last_state.s_tracking_setup .is_wysiwyg = "true";
defparam \last_state.s_tracking_setup .power_up = "low";

dffeas \last_state.s_phy_initialise (
	.clk(clk),
	.d(\state.s_phy_initialise~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_phy_initialise~q ),
	.prn(vcc));
defparam \last_state.s_phy_initialise .is_wysiwyg = "true";
defparam \last_state.s_phy_initialise .power_up = "low";

cycloneiii_lcell_comb \WideNor1~13 (
	.dataa(last_states_read_mtp),
	.datab(\last_state.s_tracking_setup~q ),
	.datac(\last_state.s_phy_initialise~q ),
	.datad(\last_state.s_tracking~q ),
	.cin(gnd),
	.combout(\WideNor1~13_combout ),
	.cout());
defparam \WideNor1~13 .lut_mask = 16'hFFFE;
defparam \WideNor1~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~14 (
	.dataa(last_states_rrp_seek),
	.datab(last_states_adv_rd_lat),
	.datac(last_states_rrp_sweep),
	.datad(\last_state.s_poa~q ),
	.cin(gnd),
	.combout(\WideNor1~14_combout ),
	.cout());
defparam \WideNor1~14 .lut_mask = 16'hFEFF;
defparam \WideNor1~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~15 (
	.dataa(last_states_adv_wr_lat),
	.datab(last_states_rrp_reset),
	.datac(\WideNor1~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideNor1~15_combout ),
	.cout());
defparam \WideNor1~15 .lut_mask = 16'hFEFE;
defparam \WideNor1~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr1~8 (
	.dataa(WideOr0),
	.datab(gnd),
	.datac(ac_muxctrl_broadcast_rcommandcmd_init_dram),
	.datad(curr_cmdcmd_prep_customer_mr_setup),
	.cin(gnd),
	.combout(\WideOr1~8_combout ),
	.cout());
defparam \WideOr1~8 .lut_mask = 16'hAFFF;
defparam \WideOr1~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideNor1~16 (
	.dataa(\WideNor1~12_combout ),
	.datab(\WideNor1~13_combout ),
	.datac(\WideNor1~15_combout ),
	.datad(\WideOr1~8_combout ),
	.cin(gnd),
	.combout(\WideNor1~16_combout ),
	.cout());
defparam \WideNor1~16 .lut_mask = 16'hFEFF;
defparam \WideNor1~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector41~0 (
	.dataa(\state.s_poa~q ),
	.datab(\WideNor1~16_combout ),
	.datac(gnd),
	.datad(\WideOr34~6_combout ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hFF77;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_5),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFFFE;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[5] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[5]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[5] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[5] .power_up = "low";

cycloneiii_lcell_comb \mtp_almt:dvw_size_a1[0]~0 (
	.dataa(\curr_ctrl.command_done~q ),
	.datab(\state.s_read_mtp~q ),
	.datac(\mtp_almts_checked[1]~q ),
	.datad(\mtp_almts_checked[0]~q ),
	.cin(gnd),
	.combout(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.cout());
defparam \mtp_almt:dvw_size_a1[0]~0 .lut_mask = 16'hFFFE;
defparam \mtp_almt:dvw_size_a1[0]~0 .sum_lutc_input = "datac";

dffeas \mtp_almt:dvw_size_a1[5] (
	.clk(clk),
	.d(\curr_ctrl.command_result[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[5]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[5] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[5] .power_up = "low";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_4),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hFFFE;
defparam \Selector5~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[4] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[4]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[4] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[4] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[4] (
	.clk(clk),
	.d(\curr_ctrl.command_result[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[4]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[4] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[4] .power_up = "low";

cycloneiii_lcell_comb \Selector6~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_3),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hFFFE;
defparam \Selector6~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[3] (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[3]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[3] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[3] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[3] (
	.clk(clk),
	.d(\curr_ctrl.command_result[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[3]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[3] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[3] .power_up = "low";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_2),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hFFFE;
defparam \Selector7~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[2] (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[2]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[2] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[2] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[2] (
	.clk(clk),
	.d(\curr_ctrl.command_result[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[2]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[2] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[2] .power_up = "low";

cycloneiii_lcell_comb \Selector8~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_1),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFFFE;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[1] (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[1]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[1] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[1] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[1] (
	.clk(clk),
	.d(\curr_ctrl.command_result[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[1]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[1] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[1] .power_up = "low";

cycloneiii_lcell_comb \Selector9~0 (
	.dataa(curr_cmdcmd_idle),
	.datab(Selector1),
	.datac(WideOr0),
	.datad(dgrb_ctrlcommand_result_0),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hFFFE;
defparam \Selector9~0 .sum_lutc_input = "datac";

dffeas \curr_ctrl.command_result[0] (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[0]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[0] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[0] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[0] (
	.clk(clk),
	.d(\curr_ctrl.command_result[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[0]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[0] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[0] .power_up = "low";

cycloneiii_lcell_comb \LessThan0~1 (
	.dataa(\mtp_almt:dvw_size_a0[0]~q ),
	.datab(\mtp_almt:dvw_size_a1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h00DD;
defparam \LessThan0~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~3 (
	.dataa(\mtp_almt:dvw_size_a0[1]~q ),
	.datab(\mtp_almt:dvw_size_a1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h00BF;
defparam \LessThan0~3 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~5 (
	.dataa(\mtp_almt:dvw_size_a0[2]~q ),
	.datab(\mtp_almt:dvw_size_a1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h00DF;
defparam \LessThan0~5 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~7 (
	.dataa(\mtp_almt:dvw_size_a0[3]~q ),
	.datab(\mtp_almt:dvw_size_a1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h00BF;
defparam \LessThan0~7 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~9 (
	.dataa(\mtp_almt:dvw_size_a0[4]~q ),
	.datab(\mtp_almt:dvw_size_a1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h00DF;
defparam \LessThan0~9 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~10 (
	.dataa(\mtp_almt:dvw_size_a0[5]~q ),
	.datab(\mtp_almt:dvw_size_a1[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~9_cout ),
	.combout(\LessThan0~10_combout ),
	.cout());
defparam \LessThan0~10 .lut_mask = 16'hFDFD;
defparam \LessThan0~10 .sum_lutc_input = "cin";

dffeas mtp_correct_almt(
	.clk(clk),
	.d(\LessThan0~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mtp_correct_almt~q ),
	.prn(vcc));
defparam mtp_correct_almt.is_wysiwyg = "true";
defparam mtp_correct_almt.power_up = "low";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_dgrb (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	clk,
	seq_ac_add_1t_ac_lat_internal,
	rst_n,
	sig_doing_rd_0,
	sig_doing_rd_1,
	dgrb_ac_access_req1,
	sig_addr_cmd0cs_n0,
	sig_addr_cmd0addr2,
	sig_addr_cmd0addr3,
	sig_addr_cmd0addr4,
	sig_addr_cmd0addr5,
	sig_addr_cmd0cas_n,
	wd_lat_0,
	wd_lat_1,
	wd_lat_4,
	wd_lat_3,
	wd_lat_2,
	dgb_ac_access_gnt_r,
	seq_rdata_valid_lat_dec1,
	seq_pll_inc_dec_n1,
	seq_pll_start_reconfig1,
	ac_muxctrl_broadcast_rcommand_req,
	dgrb_ctrlcommand_done,
	curr_cmdcmd_idle,
	WideOr1,
	last_states_rdv,
	last_states_read_mtp,
	last_states_rrp_seek,
	last_states_adv_rd_lat,
	last_states_rrp_sweep,
	last_states_adv_wr_lat,
	last_states_rrp_reset,
	rdata_valid,
	seq_pll_select_2,
	seq_pll_select_0,
	\ctrl_dgrb.command_op.single_bit ,
	\ctrl_dgrb.command_op.mtp_almt ,
	Selector57,
	Selector52,
	phs_shft_busy,
	dgrb_ctrlcommand_result_5,
	dgrb_ctrlcommand_result_4,
	dgrb_ctrlcommand_result_3,
	dgrb_ctrlcommand_result_2,
	dgrb_ctrlcommand_result_1,
	dgrb_ctrlcommand_result_0,
	mmc_seq_done,
	seq_mmc_start1,
	mimic_value_captured,
	GND_port)/* synthesis synthesis_greybox=1 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	clk;
input 	seq_ac_add_1t_ac_lat_internal;
input 	rst_n;
output 	sig_doing_rd_0;
output 	sig_doing_rd_1;
output 	dgrb_ac_access_req1;
output 	sig_addr_cmd0cs_n0;
output 	sig_addr_cmd0addr2;
output 	sig_addr_cmd0addr3;
output 	sig_addr_cmd0addr4;
output 	sig_addr_cmd0addr5;
output 	sig_addr_cmd0cas_n;
output 	wd_lat_0;
output 	wd_lat_1;
output 	wd_lat_4;
output 	wd_lat_3;
output 	wd_lat_2;
input 	dgb_ac_access_gnt_r;
output 	seq_rdata_valid_lat_dec1;
output 	seq_pll_inc_dec_n1;
output 	seq_pll_start_reconfig1;
input 	ac_muxctrl_broadcast_rcommand_req;
output 	dgrb_ctrlcommand_done;
input 	curr_cmdcmd_idle;
input 	WideOr1;
input 	last_states_rdv;
input 	last_states_read_mtp;
input 	last_states_rrp_seek;
input 	last_states_adv_rd_lat;
input 	last_states_rrp_sweep;
input 	last_states_adv_wr_lat;
input 	last_states_rrp_reset;
input 	[0:0] rdata_valid;
output 	seq_pll_select_2;
output 	seq_pll_select_0;
input 	\ctrl_dgrb.command_op.single_bit ;
input 	\ctrl_dgrb.command_op.mtp_almt ;
input 	Selector57;
input 	Selector52;
input 	phs_shft_busy;
output 	dgrb_ctrlcommand_result_5;
output 	dgrb_ctrlcommand_result_4;
output 	dgrb_ctrlcommand_result_3;
output 	dgrb_ctrlcommand_result_2;
output 	dgrb_ctrlcommand_result_1;
output 	dgrb_ctrlcommand_result_0;
input 	mmc_seq_done;
output 	seq_mmc_start1;
input 	mimic_value_captured;
input 	GND_port;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \ac_block:sig_doing_rd_count~q ;
wire \Add23~0_combout ;
wire \Add23~2_combout ;
wire \Add23~4_combout ;
wire \Add23~13 ;
wire \Add23~14_combout ;
wire \sig_trk_ack~q ;
wire \trk_block:sig_req_rsc_shift[5]~q ;
wire \trk_block:sig_req_rsc_shift[4]~q ;
wire \trk_block:sig_mimic_delta[0]~q ;
wire \Add15~0_combout ;
wire \trk_block:sig_large_drift_seen~q ;
wire \trk_block:sig_mimic_delta[5]~q ;
wire \trk_block:sig_mimic_delta[4]~q ;
wire \trk_block:sig_mimic_delta[3]~q ;
wire \trk_block:sig_mimic_delta[2]~q ;
wire \trk_block:sig_mimic_delta[1]~q ;
wire \Add15~7 ;
wire \Add15~9 ;
wire \Add15~8_combout ;
wire \Add15~11 ;
wire \Add15~10_combout ;
wire \Add15~13 ;
wire \Add15~12_combout ;
wire \Add16~2_combout ;
wire \Add16~4_combout ;
wire \Add16~6_combout ;
wire \Add16~8_combout ;
wire \Add16~10_combout ;
wire \Add16~12_combout ;
wire \Add18~7 ;
wire \Add18~9 ;
wire \Add18~8_combout ;
wire \Add18~11 ;
wire \Add18~10_combout ;
wire \Add18~13 ;
wire \Add18~12_combout ;
wire \trk_block:sig_req_rsc_shift[5]~0_combout ;
wire \trk_block:sig_req_rsc_shift[4]~0_combout ;
wire \Add15~14_combout ;
wire \Add18~14_combout ;
wire \trk_block:trk_proc:v_remaining_samples[3]~q ;
wire \trk_block:sig_rsc_drift[6]~q ;
wire \trk_block:sig_rsc_drift[5]~q ;
wire \trk_block:sig_rsc_drift[4]~q ;
wire \trk_block:sig_rsc_drift[3]~q ;
wire \trk_block:sig_rsc_drift[2]~q ;
wire \trk_block:sig_rsc_drift[1]~q ;
wire \Add9~1 ;
wire \Add9~3 ;
wire \Add9~2_combout ;
wire \Add9~5 ;
wire \Add9~4_combout ;
wire \Add9~7 ;
wire \Add9~6_combout ;
wire \Add9~9 ;
wire \Add9~8_combout ;
wire \Add9~11 ;
wire \Add9~10_combout ;
wire \Add9~13_cout ;
wire \Add9~15_cout ;
wire \Add9~16_combout ;
wire \rsc_block:sig_test_dq_expired~q ;
wire \Add5~18 ;
wire \Add5~19_combout ;
wire \Add6~1 ;
wire \Add6~3 ;
wire \Add6~2_combout ;
wire \Add6~5 ;
wire \Add6~4_combout ;
wire \Add6~7 ;
wire \Add6~6_combout ;
wire \Add6~9 ;
wire \Add6~8_combout ;
wire \Add6~11 ;
wire \Add6~10_combout ;
wire \Add6~13 ;
wire \Add6~12_combout ;
wire \Add6~14_combout ;
wire \sig_cdvw_state.current_bit[0]~q ;
wire \Add11~13 ;
wire \Add11~12_combout ;
wire \Add12~1 ;
wire \Add12~0_combout ;
wire \Add12~3 ;
wire \Add12~2_combout ;
wire \Add12~5 ;
wire \Add12~4_combout ;
wire \Add12~7 ;
wire \Add12~6_combout ;
wire \Add12~9 ;
wire \Add12~8_combout ;
wire \Add12~11 ;
wire \Add12~10_combout ;
wire \Add12~12_combout ;
wire \Add11~16 ;
wire \Add11~15_combout ;
wire \Add11~18 ;
wire \Add11~17_combout ;
wire \Add11~20 ;
wire \Add11~19_combout ;
wire \Add11~22 ;
wire \Add11~21_combout ;
wire \Add11~24 ;
wire \Add11~23_combout ;
wire \Add11~25_combout ;
wire \Add10~1 ;
wire \Add10~0_combout ;
wire \Add10~3 ;
wire \Add10~2_combout ;
wire \Add10~5 ;
wire \Add10~4_combout ;
wire \Add10~7 ;
wire \Add10~6_combout ;
wire \Add10~9 ;
wire \Add10~8_combout ;
wire \Add10~11 ;
wire \Add10~10_combout ;
wire \Add10~13 ;
wire \Add10~12_combout ;
wire \Add10~14_combout ;
wire \trk_block:trk_proc:v_remaining_samples[3]~0_combout ;
wire \Add17~3_cout ;
wire \Add17~5 ;
wire \Add17~4_combout ;
wire \Add17~7 ;
wire \Add17~6_combout ;
wire \Add17~9 ;
wire \Add17~8_combout ;
wire \Add17~11 ;
wire \Add17~10_combout ;
wire \Add17~13 ;
wire \Add17~12_combout ;
wire \Add17~15 ;
wire \Add17~14_combout ;
wire \Add17~16_combout ;
wire \trk_block:sig_rsc_drift[6]~0_combout ;
wire \trk_block:sig_rsc_drift[5]~0_combout ;
wire \trk_block:sig_rsc_drift[4]~0_combout ;
wire \trk_block:sig_rsc_drift[3]~0_combout ;
wire \trk_block:sig_rsc_drift[2]~0_combout ;
wire \trk_block:sig_rsc_drift[1]~0_combout ;
wire \sig_cdvw_state.current_window_centre[5]~q ;
wire \sig_cdvw_state.current_window_centre[4]~q ;
wire \sig_cdvw_state.current_window_centre[3]~q ;
wire \sig_cdvw_state.current_window_centre[2]~q ;
wire \sig_cdvw_state.current_window_centre[1]~q ;
wire \sig_cdvw_state.current_window_centre[0]~q ;
wire \sig_cdvw_state.current_bit[0]~6_combout ;
wire \sig_cdvw_state.current_window_centre[0]~7 ;
wire \sig_cdvw_state.current_window_centre[0]~6_combout ;
wire \sig_cdvw_state.current_window_centre[1]~9 ;
wire \sig_cdvw_state.current_window_centre[1]~8_combout ;
wire \sig_cdvw_state.current_window_centre[2]~11 ;
wire \sig_cdvw_state.current_window_centre[2]~10_combout ;
wire \sig_cdvw_state.current_window_centre[3]~13 ;
wire \sig_cdvw_state.current_window_centre[3]~12_combout ;
wire \sig_cdvw_state.current_window_centre[4]~15 ;
wire \sig_cdvw_state.current_window_centre[4]~14_combout ;
wire \sig_cdvw_state.current_window_centre[5]~16_combout ;
wire \sig_rsc_cdvw_phase~q ;
wire \ac_block:sig_count[7]~q ;
wire \Selector140~6_combout ;
wire \sig_addr_cmd[0].addr[12]~0_combout ;
wire \sig_addr_cmd[0].addr[12]~1_combout ;
wire \ac_block:sig_count[7]~3_combout ;
wire \Selector166~0_combout ;
wire \ac_block:sig_count[7]~6_combout ;
wire \Selector170~0_combout ;
wire \sig_ac_req.s_ac_read_wd_lat~q ;
wire \WideOr26~0_combout ;
wire \ac_block:sig_count[5]~1_combout ;
wire \Selector169~2_combout ;
wire \Selector169~3_combout ;
wire \Selector169~4_combout ;
wire \sig_doing_rd_count~10_combout ;
wire \Selector25~0_combout ;
wire \sig_dgrb_state.s_poa_cal~q ;
wire \Selector26~0_combout ;
wire \Selector21~0_combout ;
wire \sig_dgrb_state~244_combout ;
wire \sig_dgrb_state~245_combout ;
wire \sig_dgrb_state~248_combout ;
wire \sig_dgrb_state~249_combout ;
wire \sig_dgrb_state~250_combout ;
wire \sig_dgrb_state~252_combout ;
wire \sig_dgrb_state~253_combout ;
wire \trk_block:sig_req_rsc_shift[6]~q ;
wire \LessThan10~0_combout ;
wire \LessThan10~2_combout ;
wire \rsc_block:sig_rewind_direction~q ;
wire \rsc_block:sig_num_phase_shifts[5]~q ;
wire \rsc_block:sig_count[7]~q ;
wire \rsc_block:sig_count[6]~q ;
wire \rsc_block:sig_count[5]~q ;
wire \rsc_block:sig_count[4]~q ;
wire \Equal7~0_combout ;
wire \rsc_block:sig_count[3]~q ;
wire \rsc_block:sig_count[2]~q ;
wire \rsc_block:sig_count[1]~q ;
wire \Equal7~1_combout ;
wire \Selector59~1_combout ;
wire \sig_dgrb_state~266_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ;
wire \ctrl_dgrb_r.command.cmd_poa~q ;
wire \sig_dgrb_state~275_combout ;
wire \sig_dgrb_state~276_combout ;
wire \trk_block:sig_trk_state.s_trk_complete~q ;
wire \Selector127~0_combout ;
wire \sig_req_rsc_shift~58_combout ;
wire \trk_block:sig_mimic_delta[7]~q ;
wire \sig_req_rsc_shift~59_combout ;
wire \sig_req_rsc_shift~61_combout ;
wire \sig_req_rsc_shift~62_combout ;
wire \sig_req_rsc_shift~63_combout ;
wire \sig_req_rsc_shift~64_combout ;
wire \sig_req_rsc_shift~65_combout ;
wire \trk_block:trk_proc:v_remaining_samples[6]~q ;
wire \trk_block:sig_rsc_drift[7]~q ;
wire \cal_codvw_phase[5]~q ;
wire \cal_codvw_phase[4]~q ;
wire \cal_codvw_phase[3]~q ;
wire \cal_codvw_phase[2]~q ;
wire \cal_codvw_phase[1]~q ;
wire \trk_block:sig_rsc_drift[0]~q ;
wire \sig_rewind_direction~1_combout ;
wire \Add5~1_combout ;
wire \Add5~2_combout ;
wire \Add5~4_combout ;
wire \Add5~5_combout ;
wire \Add5~6_combout ;
wire \Add5~7_combout ;
wire \Add5~21_combout ;
wire \Selector48~0_combout ;
wire \Selector57~0_combout ;
wire \rsc_block:sig_count[6]~0_combout ;
wire \rsc_block:sig_count[6]~2_combout ;
wire \Selector39~0_combout ;
wire \rsc_block:sig_count[6]~3_combout ;
wire \rsc_block:sig_count[6]~4_combout ;
wire \Selector40~0_combout ;
wire \sig_cdvw_state.largest_window_centre[5]~q ;
wire \Selector41~0_combout ;
wire \Selector42~2_combout ;
wire \sig_cdvw_state.largest_window_centre[4]~q ;
wire \Selector43~0_combout ;
wire \sig_cdvw_state.largest_window_centre[3]~q ;
wire \Selector43~1_combout ;
wire \Selector43~2_combout ;
wire \Selector44~0_combout ;
wire \sig_cdvw_state.largest_window_centre[2]~q ;
wire \Selector44~1_combout ;
wire \Selector45~0_combout ;
wire \sig_cdvw_state.largest_window_centre[1]~q ;
wire \Selector45~1_combout ;
wire \Selector56~0_combout ;
wire \find_centre_of_largest_data_valid_window~5_combout ;
wire \find_centre_of_largest_data_valid_window~0_combout ;
wire \sig_cdvw_state.first_good_edge[2]~q ;
wire \sig_cdvw_state.first_good_edge[5]~q ;
wire \v_cdvw_state~424_combout ;
wire \sig_cdvw_state.invalid_phase_seen~q ;
wire \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ;
wire \Selector51~2_combout ;
wire \sig_trk_state~116_combout ;
wire \sig_trk_state~120_combout ;
wire \trk_block:sig_mimic_cdv[0]~q ;
wire \Add11~14_combout ;
wire \trk_proc~6_combout ;
wire \LessThan7~0_combout ;
wire \LessThan7~1_combout ;
wire \trk_block:sig_mimic_cdv[5]~q ;
wire \trk_block:sig_mimic_cdv[4]~q ;
wire \trk_block:sig_mimic_cdv[3]~q ;
wire \trk_block:sig_mimic_cdv[2]~q ;
wire \trk_block:sig_mimic_cdv[1]~q ;
wire \Add11~27_combout ;
wire \Selector119~0_combout ;
wire \Selector119~1_combout ;
wire \Selector119~2_combout ;
wire \Selector122~0_combout ;
wire \Add17~18_combout ;
wire \Add17~19_combout ;
wire \Add17~20_combout ;
wire \Selector95~0_combout ;
wire \Add17~21_combout ;
wire \sig_rsc_drift~40_combout ;
wire \Selector96~0_combout ;
wire \Add17~22_combout ;
wire \sig_rsc_drift~41_combout ;
wire \Selector69~2_combout ;
wire \Selector97~0_combout ;
wire \Add17~23_combout ;
wire \sig_rsc_drift~42_combout ;
wire \Selector70~0_combout ;
wire \Selector98~0_combout ;
wire \Add17~24_combout ;
wire \sig_rsc_drift~43_combout ;
wire \Selector71~0_combout ;
wire \Selector99~0_combout ;
wire \Add17~25_combout ;
wire \sig_rsc_drift~44_combout ;
wire \Selector72~0_combout ;
wire \Selector100~0_combout ;
wire \Add17~26_combout ;
wire \sig_rsc_drift~45_combout ;
wire \Selector73~0_combout ;
wire \Add17~27_combout ;
wire \sig_test_dq_expired~6_combout ;
wire \Equal8~0_combout ;
wire \v_cdvw_state~434_combout ;
wire \v_cdvw_state~435_combout ;
wire \v_cdvw_state~436_combout ;
wire \v_cdvw_state~437_combout ;
wire \v_cdvw_state~438_combout ;
wire \v_cdvw_state~441_combout ;
wire \v_cdvw_state~442_combout ;
wire \v_cdvw_state~447_combout ;
wire \v_cdvw_state~450_combout ;
wire \Selector50~0_combout ;
wire \tp_match_block:sig_rdata_valid_2t~q ;
wire \trk_block:sig_mimic_cdv[0]~1_combout ;
wire \Selector35~0_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \sig_cdvw_state.current_window_centre[5]~18_combout ;
wire \sig_cdvw_state.current_window_centre[5]~19_combout ;
wire \sig_cdvw_state.current_window_centre[5]~20_combout ;
wire \sig_cdvw_state.window_centre_update~q ;
wire \sig_cdvw_state.current_window_centre[5]~21_combout ;
wire \sig_cdvw_state.current_window_centre[5]~22_combout ;
wire \sig_cdvw_state.current_window_size[0]~19_combout ;
wire \v_cdvw_state~464_combout ;
wire \v_cdvw_state~465_combout ;
wire \trk_block:sig_trk_last_state.s_trk_mimic_sample~q ;
wire \sig_trk_last_state~31_combout ;
wire \sig_trk_cdvw_phase~q ;
wire \v_cdvw_state~528_combout ;
wire \v_cdvw_state~529_combout ;
wire \sig_trk_cdvw_phase~1_combout ;
wire \rsc_block:rsc_proc:v_phase_works~q ;
wire \rsc_proc~3_combout ;
wire \sig_rsc_cdvw_phase~5_combout ;
wire \Selector66~0_combout ;
wire \Selector66~1_combout ;
wire \sig_req_rsc_shift~68_combout ;
wire \Selector42~3_combout ;
wire \Add11~28_combout ;
wire \Add11~29_combout ;
wire \Add11~30_combout ;
wire \Add11~31_combout ;
wire \Add11~32_combout ;
wire \Add11~33_combout ;
wire \Add23~1 ;
wire \Add23~3 ;
wire \Add23~5 ;
wire \Add23~7 ;
wire \Add23~9 ;
wire \Add23~11 ;
wire \Add23~12_combout ;
wire \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ;
wire \sig_dgrb_state~237_combout ;
wire \sig_dgrb_state~261_combout ;
wire \sig_dgrb_state~262_combout ;
wire \sig_dgrb_state~264_combout ;
wire \sig_dgrb_state~281_combout ;
wire \sig_dgrb_state.s_adv_wd_lat~q ;
wire \sig_dgrb_state~268_combout ;
wire \sig_dgrb_state~269_combout ;
wire \sig_dgrb_state~259_combout ;
wire \sig_dgrb_state.s_reset_cdvw~q ;
wire \sig_rsc_req~28_combout ;
wire \sig_rsc_req.s_rsc_reset_cdvw~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_idle~q ;
wire \Selector54~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ;
wire \Selector37~0_combout ;
wire \WideOr12~0_combout ;
wire \sig_dq_pin_ctr[3]~16_combout ;
wire \sig_dq_pin_ctr[1]~q ;
wire \Equal4~2_combout ;
wire \Selector36~0_combout ;
wire \sig_dq_pin_ctr[2]~q ;
wire \Equal4~1_combout ;
wire \Selector35~1_combout ;
wire \sig_dq_pin_ctr[3]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \Mux0~9_combout ;
wire \tp_match_block:sig_rdata_current_pin[14]~q ;
wire \tp_match_block:sig_rdata_current_pin[13]~q ;
wire \tp_match_block:sig_rdata_current_pin[11]~q ;
wire \tp_match_block:sig_rdata_current_pin[9]~q ;
wire \tp_match_block:sig_rdata_current_pin[12]~q ;
wire \tp_match_block:sig_rdata_current_pin[10]~q ;
wire \tp_match_block:sig_rdata_current_pin[8]~q ;
wire \Equal8~1_combout ;
wire \tp_match_block:sig_rdata_current_pin[6]~q ;
wire \tp_match_block:sig_rdata_current_pin[7]~q ;
wire \tp_match_block:sig_rdata_current_pin[5]~q ;
wire \tp_match_block:sig_rdata_current_pin[4]~q ;
wire \Equal8~2_combout ;
wire \tp_match_block:sig_rdata_current_pin[2]~q ;
wire \tp_match_block:sig_rdata_current_pin[0]~q ;
wire \tp_match_block:sig_rdata_current_pin[3]~q ;
wire \tp_match_block:sig_rdata_current_pin[1]~q ;
wire \Equal8~3_combout ;
wire \Equal8~4_combout ;
wire \sig_mtp_match~q ;
wire \rsc_block:sig_curr_byte_ln_dis~q ;
wire \rsc_proc~1_combout ;
wire \Selector51~0_combout ;
wire \Selector52~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_test_dq~q ;
wire \rsc_block:sig_num_phase_shifts[2]~0_combout ;
wire \Equal4~0_combout ;
wire \rsc_block:sig_chkd_all_dq_pins~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ;
wire \Selector51~1_combout ;
wire \Selector48~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_next_phase~q ;
wire \Add5~3_combout ;
wire \Add5~9_combout ;
wire \Add5~26_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~1_combout ;
wire \phs_shft_busy_reg:phs_shft_busy_1r~q ;
wire \phs_shft_busy_reg:phs_shft_busy_2r~q ;
wire \sig_phs_shft_busy~q ;
wire \sig_phs_shft_busy_1t~q ;
wire \rsc_block:sig_num_phase_shifts[2]~2_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~3_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~4_combout ;
wire \rsc_block:sig_num_phase_shifts[0]~q ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ;
wire \trk_block:sig_mmc_seq_done_1t~q ;
wire \trk_block:trk_proc:v_remaining_samples[2]~0_combout ;
wire \ctrl_dgrb_r.command.cmd_tr_due~q ;
wire \sig_dgrb_state~241_combout ;
wire \sig_dgrb_state.s_track~q ;
wire \sig_dgrb_last_state.s_track~q ;
wire \cdvw_proc~1_combout ;
wire \v_cdvw_state~430_combout ;
wire \v_cdvw_state~461_combout ;
wire \sig_cdvw_state.largest_window_size[0]~1_combout ;
wire \sig_cdvw_state.largest_window_size[1]~q ;
wire \sig_cdvw_state.current_window_size[0]~7 ;
wire \sig_cdvw_state.current_window_size[1]~8_combout ;
wire \cdvw_proc~2_combout ;
wire \v_cdvw_state~530_combout ;
wire \sig_rsc_cdvw_shift_in~4_combout ;
wire \sig_rsc_cdvw_shift_in~q ;
wire \shift_in_mmc_seq_value~0_combout ;
wire \sig_trk_cdvw_shift_in~q ;
wire \sig_cdvw_state.working_window[12]~4_combout ;
wire \sig_cdvw_state.working_window[12]~5_combout ;
wire \v_cdvw_state~531_combout ;
wire \sig_cdvw_state.working_window[63]~q ;
wire \v_cdvw_state~527_combout ;
wire \sig_cdvw_state.working_window[12]~6_combout ;
wire \sig_cdvw_state.working_window[62]~q ;
wire \v_cdvw_state~526_combout ;
wire \sig_cdvw_state.working_window[61]~q ;
wire \v_cdvw_state~525_combout ;
wire \sig_cdvw_state.working_window[60]~q ;
wire \v_cdvw_state~524_combout ;
wire \sig_cdvw_state.working_window[59]~q ;
wire \v_cdvw_state~523_combout ;
wire \sig_cdvw_state.working_window[58]~q ;
wire \v_cdvw_state~522_combout ;
wire \sig_cdvw_state.working_window[57]~q ;
wire \v_cdvw_state~521_combout ;
wire \sig_cdvw_state.working_window[56]~q ;
wire \v_cdvw_state~520_combout ;
wire \sig_cdvw_state.working_window[55]~q ;
wire \v_cdvw_state~519_combout ;
wire \sig_cdvw_state.working_window[54]~q ;
wire \v_cdvw_state~518_combout ;
wire \sig_cdvw_state.working_window[53]~q ;
wire \v_cdvw_state~517_combout ;
wire \sig_cdvw_state.working_window[52]~q ;
wire \v_cdvw_state~516_combout ;
wire \sig_cdvw_state.working_window[51]~q ;
wire \v_cdvw_state~515_combout ;
wire \sig_cdvw_state.working_window[50]~q ;
wire \v_cdvw_state~514_combout ;
wire \sig_cdvw_state.working_window[49]~q ;
wire \v_cdvw_state~513_combout ;
wire \sig_cdvw_state.working_window[48]~q ;
wire \v_cdvw_state~512_combout ;
wire \sig_cdvw_state.working_window[47]~q ;
wire \v_cdvw_state~511_combout ;
wire \sig_cdvw_state.working_window[46]~q ;
wire \v_cdvw_state~510_combout ;
wire \sig_cdvw_state.working_window[45]~q ;
wire \v_cdvw_state~509_combout ;
wire \sig_cdvw_state.working_window[44]~q ;
wire \v_cdvw_state~508_combout ;
wire \sig_cdvw_state.working_window[43]~q ;
wire \v_cdvw_state~507_combout ;
wire \sig_cdvw_state.working_window[42]~q ;
wire \v_cdvw_state~506_combout ;
wire \sig_cdvw_state.working_window[41]~q ;
wire \v_cdvw_state~505_combout ;
wire \sig_cdvw_state.working_window[40]~q ;
wire \v_cdvw_state~504_combout ;
wire \sig_cdvw_state.working_window[39]~q ;
wire \v_cdvw_state~503_combout ;
wire \sig_cdvw_state.working_window[38]~q ;
wire \v_cdvw_state~502_combout ;
wire \sig_cdvw_state.working_window[37]~q ;
wire \v_cdvw_state~501_combout ;
wire \sig_cdvw_state.working_window[36]~q ;
wire \v_cdvw_state~500_combout ;
wire \sig_cdvw_state.working_window[35]~q ;
wire \v_cdvw_state~499_combout ;
wire \sig_cdvw_state.working_window[34]~q ;
wire \v_cdvw_state~498_combout ;
wire \sig_cdvw_state.working_window[33]~q ;
wire \v_cdvw_state~497_combout ;
wire \sig_cdvw_state.working_window[32]~q ;
wire \v_cdvw_state~496_combout ;
wire \sig_cdvw_state.working_window[31]~q ;
wire \v_cdvw_state~495_combout ;
wire \sig_cdvw_state.working_window[30]~q ;
wire \v_cdvw_state~494_combout ;
wire \sig_cdvw_state.working_window[29]~q ;
wire \v_cdvw_state~493_combout ;
wire \sig_cdvw_state.working_window[28]~q ;
wire \v_cdvw_state~492_combout ;
wire \sig_cdvw_state.working_window[27]~q ;
wire \v_cdvw_state~491_combout ;
wire \sig_cdvw_state.working_window[26]~q ;
wire \v_cdvw_state~490_combout ;
wire \sig_cdvw_state.working_window[25]~q ;
wire \v_cdvw_state~489_combout ;
wire \sig_cdvw_state.working_window[24]~q ;
wire \v_cdvw_state~488_combout ;
wire \sig_cdvw_state.working_window[23]~q ;
wire \v_cdvw_state~487_combout ;
wire \sig_cdvw_state.working_window[22]~q ;
wire \v_cdvw_state~486_combout ;
wire \sig_cdvw_state.working_window[21]~q ;
wire \v_cdvw_state~485_combout ;
wire \sig_cdvw_state.working_window[20]~q ;
wire \v_cdvw_state~484_combout ;
wire \sig_cdvw_state.working_window[19]~q ;
wire \v_cdvw_state~483_combout ;
wire \sig_cdvw_state.working_window[18]~q ;
wire \v_cdvw_state~482_combout ;
wire \sig_cdvw_state.working_window[17]~q ;
wire \v_cdvw_state~481_combout ;
wire \sig_cdvw_state.working_window[16]~q ;
wire \v_cdvw_state~480_combout ;
wire \sig_cdvw_state.working_window[15]~q ;
wire \v_cdvw_state~479_combout ;
wire \sig_cdvw_state.working_window[14]~q ;
wire \v_cdvw_state~478_combout ;
wire \sig_cdvw_state.working_window[13]~q ;
wire \v_cdvw_state~477_combout ;
wire \sig_cdvw_state.working_window[12]~q ;
wire \v_cdvw_state~476_combout ;
wire \sig_cdvw_state.working_window[11]~q ;
wire \v_cdvw_state~475_combout ;
wire \sig_cdvw_state.working_window[10]~q ;
wire \v_cdvw_state~474_combout ;
wire \sig_cdvw_state.working_window[9]~q ;
wire \v_cdvw_state~473_combout ;
wire \sig_cdvw_state.working_window[8]~q ;
wire \v_cdvw_state~472_combout ;
wire \sig_cdvw_state.working_window[7]~q ;
wire \v_cdvw_state~471_combout ;
wire \sig_cdvw_state.working_window[6]~q ;
wire \v_cdvw_state~470_combout ;
wire \sig_cdvw_state.working_window[5]~q ;
wire \v_cdvw_state~469_combout ;
wire \sig_cdvw_state.working_window[4]~q ;
wire \v_cdvw_state~468_combout ;
wire \sig_cdvw_state.working_window[3]~q ;
wire \v_cdvw_state~467_combout ;
wire \sig_cdvw_state.working_window[2]~q ;
wire \v_cdvw_state~466_combout ;
wire \sig_cdvw_state.working_window[1]~q ;
wire \v_cdvw_state~463_combout ;
wire \sig_cdvw_state.working_window[0]~q ;
wire \v_cdvw_state~456_combout ;
wire \sig_cdvw_state.last_bit_value~q ;
wire \find_centre_of_largest_data_valid_window~7_combout ;
wire \sig_cdvw_state.current_window_size[0]~18_combout ;
wire \sig_cdvw_state.current_window_size[0]~20_combout ;
wire \sig_cdvw_state.current_window_size[1]~q ;
wire \sig_cdvw_state.current_window_size[1]~9 ;
wire \sig_cdvw_state.current_window_size[2]~11 ;
wire \sig_cdvw_state.current_window_size[3]~12_combout ;
wire \sig_cdvw_state.current_window_size[3]~q ;
wire \v_cdvw_state~451_combout ;
wire \v_cdvw_state~462_combout ;
wire \sig_cdvw_state.largest_window_size[0]~q ;
wire \sig_cdvw_state.current_window_size[0]~6_combout ;
wire \sig_cdvw_state.current_window_size[0]~q ;
wire \sig_cdvw_state.current_window_size[3]~13 ;
wire \sig_cdvw_state.current_window_size[4]~14_combout ;
wire \sig_cdvw_state.current_window_size[4]~q ;
wire \v_cdvw_state~452_combout ;
wire \sig_cdvw_state.current_window_size[4]~15 ;
wire \sig_cdvw_state.current_window_size[5]~16_combout ;
wire \sig_cdvw_state.current_window_size[5]~q ;
wire \sig_cdvw_state.current_window_size[2]~10_combout ;
wire \sig_cdvw_state.current_window_size[2]~q ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~10_combout ;
wire \v_cdvw_state~453_combout ;
wire \v_cdvw_state~454_combout ;
wire \v_cdvw_state~443_combout ;
wire \find_centre_of_largest_data_valid_window~6_combout ;
wire \v_cdvw_state~440_combout ;
wire \sig_cdvw_state.found_a_good_edge~q ;
wire \sig_cdvw_state.first_good_edge[1]~0_combout ;
wire \sig_cdvw_state.first_good_edge[0]~q ;
wire \sig_cdvw_state.current_bit[0]~7 ;
wire \sig_cdvw_state.current_bit[1]~11_combout ;
wire \sig_cdvw_state.current_bit[1]~12 ;
wire \sig_cdvw_state.current_bit[2]~13_combout ;
wire \sig_cdvw_state.current_bit[5]~10_combout ;
wire \sig_cdvw_state.current_bit[2]~q ;
wire \sig_cdvw_state.current_bit[2]~14 ;
wire \sig_cdvw_state.current_bit[3]~15_combout ;
wire \sig_cdvw_state.current_bit[3]~q ;
wire \sig_cdvw_state.current_bit[5]~8_combout ;
wire \sig_cdvw_state.current_bit[3]~16 ;
wire \sig_cdvw_state.current_bit[4]~17_combout ;
wire \sig_cdvw_state.current_bit[4]~q ;
wire \sig_cdvw_state.current_bit[4]~18 ;
wire \sig_cdvw_state.current_bit[5]~19_combout ;
wire \sig_cdvw_state.current_bit[5]~q ;
wire \sig_cdvw_state.current_bit[5]~9_combout ;
wire \sig_cdvw_state.current_bit[1]~q ;
wire \v_cdvw_state~444_combout ;
wire \sig_cdvw_state.first_good_edge[1]~q ;
wire \v_cdvw_state~425_combout ;
wire \v_cdvw_state~445_combout ;
wire \sig_cdvw_state.first_good_edge[3]~q ;
wire \v_cdvw_state~446_combout ;
wire \sig_cdvw_state.first_good_edge[4]~q ;
wire \v_cdvw_state~426_combout ;
wire \v_cdvw_state~427_combout ;
wire \v_cdvw_state~448_combout ;
wire \sig_cdvw_state.valid_phase_seen~q ;
wire \v_cdvw_state~428_combout ;
wire \v_cdvw_state~449_combout ;
wire \sig_cdvw_state.first_cycle~q ;
wire \v_cdvw_state~429_combout ;
wire \v_cdvw_state~433_combout ;
wire \sig_cdvw_state.status.calculating~q ;
wire \sig_cdvw_state.largest_window_size[0]~0_combout ;
wire \v_cdvw_state~455_combout ;
wire \sig_cdvw_state.multiple_eq_windows~q ;
wire \v_cdvw_state~431_combout ;
wire \v_cdvw_state~432_combout ;
wire \sig_cdvw_state.status.valid_result~q ;
wire \sig_trk_state~127_combout ;
wire \trk_block:sig_trk_state.s_trk_idle~q ;
wire \Selector123~0_combout ;
wire \Selector86~0_combout ;
wire \sig_trk_state~128_combout ;
wire \sig_trk_state~121_combout ;
wire \sig_trk_state~122_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_wait~q ;
wire \sig_phs_shft_end~0_combout ;
wire \sig_phs_shft_end~q ;
wire \sig_trk_state~109_combout ;
wire \sig_trk_last_state~29_combout ;
wire \trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ;
wire \sig_trk_state~107_combout ;
wire \sig_trk_state~114_combout ;
wire \trk_block:sig_trk_state.s_trk_adjust_resync~q ;
wire \sig_trk_state~108_combout ;
wire \sig_trk_last_state~30_combout ;
wire \trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ;
wire \sig_trk_state~110_combout ;
wire \sig_trk_state~117_combout ;
wire \sig_trk_state~118_combout ;
wire \Selector127~1_combout ;
wire \sig_trk_state~119_combout ;
wire \Selector93~0_combout ;
wire \trk_block:sig_mimic_cdv[0]~0_combout ;
wire \Selector93~1_combout ;
wire \trk_block:sig_mimic_cdv_found~q ;
wire \sig_trk_state~123_combout ;
wire \sig_trk_state~124_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_drift~q ;
wire \sig_trk_state~111_combout ;
wire \sig_trk_state~112_combout ;
wire \sig_trk_state~113_combout ;
wire \sig_trk_state~115_combout ;
wire \trk_block:sig_trk_state.s_trk_next_phase~q ;
wire \Selector86~1_combout ;
wire \trk_block:sig_trk_state.s_trk_mimic_sample~q ;
wire \trk_block:trk_proc:v_remaining_samples[2]~q ;
wire \trk_block:trk_proc:v_remaining_samples[1]~0_combout ;
wire \Selector124~0_combout ;
wire \trk_block:trk_proc:v_remaining_samples[1]~q ;
wire \trk_block:trk_proc:v_remaining_samples[0]~0_combout ;
wire \Selector125~0_combout ;
wire \trk_block:trk_proc:v_remaining_samples[0]~q ;
wire \Equal10~1_combout ;
wire \v_remaining_samples~18_combout ;
wire \trk_block:trk_proc:v_remaining_samples[7]~0_combout ;
wire \Selector118~0_combout ;
wire \trk_block:trk_proc:v_remaining_samples[7]~q ;
wire \trk_block:trk_proc:v_remaining_samples[5]~0_combout ;
wire \Selector120~0_combout ;
wire \trk_block:trk_proc:v_remaining_samples[5]~q ;
wire \trk_block:trk_proc:v_remaining_samples[4]~0_combout ;
wire \Selector121~0_combout ;
wire \trk_block:trk_proc:v_remaining_samples[4]~q ;
wire \Equal10~0_combout ;
wire \sig_trk_state~125_combout ;
wire \sig_trk_state~126_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_calc~q ;
wire \sig_trk_cdvw_calc~4_combout ;
wire \sig_trk_cdvw_calc~q ;
wire \sig_dgrb_state~258_combout ;
wire \sig_dgrb_state.s_seek_cdvw~q ;
wire \sig_dgrb_state~274_combout ;
wire \sig_dgrb_state.s_read_mtp~q ;
wire \sig_rsc_req~29_combout ;
wire \sig_rsc_req.s_rsc_cdvw_calc~q ;
wire \Selector55~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ;
wire \Selector55~1_combout ;
wire \sig_rsc_cdvw_calc~q ;
wire \sig_dgrb_state~260_combout ;
wire \sig_dgrb_state.s_test_phases~q ;
wire \WideOr11~2_combout ;
wire \Selector32~0_combout ;
wire \cdvw_block:sig_cdvw_calc_1t~q ;
wire \v_cdvw_state~439_combout ;
wire \sig_cdvw_state.largest_window_centre[0]~q ;
wire \Selector74~0_combout ;
wire \Add6~0_combout ;
wire \rsc_block:sig_count[6]~1_combout ;
wire \rsc_block:sig_count[5]~1_combout ;
wire \rsc_block:sig_count[5]~2_combout ;
wire \Selector46~0_combout ;
wire \rsc_block:sig_count[6]~5_combout ;
wire \rsc_block:sig_count[5]~3_combout ;
wire \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ;
wire \Selector69~0_combout ;
wire \WideOr13~1_combout ;
wire \rsc_block:sig_count[5]~0_combout ;
wire \rsc_block:sig_count[5]~4_combout ;
wire \rsc_block:sig_count[0]~q ;
wire \Equal7~2_combout ;
wire \Selector57~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ;
wire \Selector69~3_combout ;
wire \cal_codvw_phase[0]~q ;
wire \Add9~0_combout ;
wire \Add5~8_combout ;
wire \Add5~10 ;
wire \Add5~11_combout ;
wire \Add5~25_combout ;
wire \rsc_block:sig_num_phase_shifts[1]~q ;
wire \Equal6~1_combout ;
wire \Selector53~0_combout ;
wire \Selector53~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ;
wire \Selector69~1_combout ;
wire \Selector83~4_combout ;
wire \Selector83~5_combout ;
wire \sig_rsc_ack~q ;
wire \Selector23~0_combout ;
wire \sig_rsc_req.s_rsc_test_phase~q ;
wire \Selector47~0_combout ;
wire \Selector47~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_idle~q ;
wire \Selector49~0_combout ;
wire \Selector49~1_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_test_phase~q ;
wire \ctrl_dgrb_r.command_op.single_bit~q ;
wire \single_bit_cal~q ;
wire \Selector38~0_combout ;
wire \sig_dq_pin_ctr[0]~q ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~9_combout ;
wire \tp_match_block:sig_rdata_current_pin[15]~q ;
wire \Equal9~0_combout ;
wire \sig_poa_match~q ;
wire \tp_match_block:sig_rdata_valid_1t~q ;
wire \poa_match_proc~0_combout ;
wire \sig_poa_match_en~q ;
wire \sig_poa_state~4_combout ;
wire \poa_block:sig_poa_state~q ;
wire \sig_poa_ack~3_combout ;
wire \sig_poa_ack~q ;
wire \sig_dgrb_state~246_combout ;
wire \sig_dgrb_state~247_combout ;
wire \sig_rsc_req~27_combout ;
wire \sig_dgrb_state~242_combout ;
wire \sig_dgrb_state~270_combout ;
wire \sig_dgrb_last_state.s_adv_wd_lat~q ;
wire \sig_dgrb_state~251_combout ;
wire \sig_dgrb_state~255_combout ;
wire \sig_dgrb_state~271_combout ;
wire \sig_dgrb_state~272_combout ;
wire \sig_dgrb_state.s_adv_rd_lat~q ;
wire \sig_dgrb_state~254_combout ;
wire \sig_dgrb_state~256_combout ;
wire \sig_dgrb_state~257_combout ;
wire \sig_dgrb_state~263_combout ;
wire \sig_dgrb_state.s_idle~q ;
wire \dgrb_state_proc~4_combout ;
wire \sig_dgrb_state~265_combout ;
wire \sig_dgrb_state.s_adv_rd_lat_setup~q ;
wire \sig_dgrb_state~243_combout ;
wire \sig_dgrb_last_state.s_adv_rd_lat_setup~q ;
wire \sig_dgrb_state~267_combout ;
wire \sig_dgrb_state~239_combout ;
wire \sig_dgrb_state~273_combout ;
wire \sig_dgrb_state.s_wait_admin~q ;
wire \sig_dgrb_state~238_combout ;
wire \sig_dgrb_state~240_combout ;
wire \sig_dgrb_state.s_rdata_valid_align~q ;
wire \sig_dgrb_state~277_combout ;
wire \sig_dgrb_state~278_combout ;
wire \sig_dgrb_state~282_combout ;
wire \sig_dgrb_state~279_combout ;
wire \sig_dgrb_state~280_combout ;
wire \sig_dgrb_state.s_release_admin~q ;
wire \Selector21~1_combout ;
wire \sig_ac_req.s_ac_idle~q ;
wire \Selector24~0_combout ;
wire \Selector25~1_combout ;
wire \Selector24~1_combout ;
wire \sig_ac_req.s_ac_read_rdv~q ;
wire \sig_addr_cmd_state~39_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ;
wire \WideOr26~1_combout ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ;
wire \Selector175~10_combout ;
wire \Selector25~2_combout ;
wire \sig_ac_req.s_ac_read_poa_mtp~q ;
wire \sig_addr_cmd_state~42_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_relax~q ;
wire \ac_block:sig_count[7]~1_combout ;
wire \ac_block:sig_count[7]~2_combout ;
wire \ac_block:sig_count[5]~2_combout ;
wire \Selector168~0_combout ;
wire \ac_block:sig_count[7]~0_combout ;
wire \Selector173~0_combout ;
wire \ac_block:sig_count[5]~0_combout ;
wire \ac_block:sig_count[5]~3_combout ;
wire \ac_block:sig_count[5]~4_combout ;
wire \ac_block:sig_count[0]~q ;
wire \sig_burst_count~4_combout ;
wire \ac_block:sig_burst_count[0]~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ;
wire \ac_block:sig_count[7]~4_combout ;
wire \ac_block:sig_count[1]~0_combout ;
wire \ac_block:sig_count[7]~7_combout ;
wire \ac_block:sig_count[1]~1_combout ;
wire \ac_block:sig_count[1]~2_combout ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ;
wire \ac_block:sig_count[7]~8_combout ;
wire \ac_block:sig_count[1]~3_combout ;
wire \ac_block:sig_count[1]~q ;
wire \Equal13~1_combout ;
wire \sig_addr_cmd_state~38_combout ;
wire \sig_addr_cmd_state~44_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_relax~q ;
wire \WideOr26~2_combout ;
wire \sig_addr_cmd_state~43_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_idle~q ;
wire \ac_block:sig_setup[0]~1_combout ;
wire \ac_block:sig_setup[0]~2 ;
wire \ac_block:sig_setup[1]~2 ;
wire \ac_block:sig_setup[2]~2 ;
wire \ac_block:sig_setup[3]~1_combout ;
wire \ac_block:sig_setup[3]~q ;
wire \ac_block:sig_setup[3]~2 ;
wire \ac_block:sig_setup[4]~2_combout ;
wire \ac_block:sig_setup[4]~q ;
wire \dimm_driving_dq_proc~1_combout ;
wire \ac_block:sig_setup[4]~1_combout ;
wire \ac_block:sig_setup[0]~q ;
wire \ac_block:sig_setup[1]~1_combout ;
wire \ac_block:sig_setup[1]~q ;
wire \ac_block:sig_setup[2]~1_combout ;
wire \ac_block:sig_setup[2]~q ;
wire \Selector128~0_combout ;
wire \Selector128~1_combout ;
wire \Selector128~2_combout ;
wire \sig_dimm_driving_dq~q ;
wire \Selector52~0_combout ;
wire \Selector51~3_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ;
wire \WideOr13~0_combout ;
wire \sig_rsc_ac_access_req~q ;
wire \Selector23~1_combout ;
wire \sig_ac_req.s_ac_read_mtp~q ;
wire \sig_addr_cmd_state~40_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ;
wire \ac_block:sig_count[7]~5_combout ;
wire \Selector167~0_combout ;
wire \ac_block:sig_count[6]~q ;
wire \Add23~6_combout ;
wire \Selector170~1_combout ;
wire \ac_block:sig_count[3]~q ;
wire \Selector171~0_combout ;
wire \ac_block:sig_count[2]~q ;
wire \Selector175~3_combout ;
wire \Selector175~4_combout ;
wire \Add23~10_combout ;
wire \Selector168~1_combout ;
wire \ac_block:sig_count[5]~q ;
wire \Add23~8_combout ;
wire \Selector169~0_combout ;
wire \sig_count~171_combout ;
wire \Selector169~1_combout ;
wire \Selector169~5_combout ;
wire \Selector169~6_combout ;
wire \Selector169~7_combout ;
wire \ac_block:sig_count[4]~q ;
wire \Selector175~5_combout ;
wire \sig_addr_cmd_state~41_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ;
wire \Selector174~0_combout ;
wire \Selector174~1_combout ;
wire \Selector174~2_combout ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ;
wire \Selector175~6_combout ;
wire \Selector175~7_combout ;
wire \Selector175~8_combout ;
wire \Selector175~9_combout ;
wire \Selector165~0_combout ;
wire \Equal13~0_combout ;
wire \Selector165~1_combout ;
wire \Selector165~2_combout ;
wire \Selector141~0_combout ;
wire \Selector141~1_combout ;
wire \Selector141~2_combout ;
wire \btp_addr_array~0_combout ;
wire \ac_block:btp_addr_array[0][4]~q ;
wire \Selector141~3_combout ;
wire \Selector141~4_combout ;
wire \Selector141~5_combout ;
wire \sig_addr_cmd~435_combout ;
wire \ctrl_dgrb_r.command_op.mtp_almt~q ;
wire \current_mtp_almt~q ;
wire \ac_block:btp_addr_array[0][3]~q ;
wire \Selector140~4_combout ;
wire \Selector140~5_combout ;
wire \Selector140~7_combout ;
wire \Selector140~8_combout ;
wire \Selector139~5_combout ;
wire \sig_addr_cmd~436_combout ;
wire \Selector139~4_combout ;
wire \Selector139~9_combout ;
wire \Selector139~6_combout ;
wire \Selector139~10_combout ;
wire \Selector139~7_combout ;
wire \Selector139~8_combout ;
wire \Selector138~1_combout ;
wire \Selector138~2_combout ;
wire \sig_addr_cmd~434_combout ;
wire \Selector140~9_combout ;
wire \Selector138~0_combout ;
wire \Selector138~3_combout ;
wire \sig_addr_cmd[0].addr[12]~2_combout ;
wire \sig_addr_cmd[0].addr[12]~3_combout ;
wire \sig_addr_cmd[0].cas_n~0_combout ;
wire \sig_wd_lat~10_combout ;
wire \dgrb_main_block:sig_wd_lat[4]~0_combout ;
wire \dgrb_main_block:sig_wd_lat[0]~q ;
wire \wd_lat[0]~0_combout ;
wire \sig_wd_lat~11_combout ;
wire \dgrb_main_block:sig_wd_lat[1]~q ;
wire \sig_wd_lat~12_combout ;
wire \dgrb_main_block:sig_wd_lat[4]~q ;
wire \sig_wd_lat~13_combout ;
wire \dgrb_main_block:sig_wd_lat[3]~q ;
wire \sig_wd_lat~14_combout ;
wire \dgrb_main_block:sig_wd_lat[2]~q ;
wire \wd_lat[2]~1_combout ;
wire \seq_rdata_valid_lat_dec~3_combout ;
wire \seq_rdata_valid_lat_dec~4_combout ;
wire \pll_reconf_mux~1_combout ;
wire \sig_trk_pll_inc_dec_n~4_combout ;
wire \trk_block:sig_trk_last_state.s_trk_adjust_resync~q ;
wire \sig_trk_pll_inc_dec_n~5_combout ;
wire \sig_trk_pll_inc_dec_n~q ;
wire \Add5~12 ;
wire \Add5~14 ;
wire \Add5~16 ;
wire \Add5~17_combout ;
wire \Add5~22_combout ;
wire \rsc_block:sig_num_phase_shifts[4]~q ;
wire \Add5~15_combout ;
wire \Add5~23_combout ;
wire \rsc_block:sig_num_phase_shifts[3]~q ;
wire \Add5~13_combout ;
wire \Add5~24_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~q ;
wire \Equal6~0_combout ;
wire \Selector59~0_combout ;
wire \sig_rsc_pll_inc_dec_n~2_combout ;
wire \sig_rsc_pll_inc_dec_n~q ;
wire \seq_pll_inc_dec_n~2_combout ;
wire \Selector59~2_combout ;
wire \sig_rsc_pll_start_reconfig~q ;
wire \Add16~1 ;
wire \Add16~3 ;
wire \Add16~5 ;
wire \Add16~7 ;
wire \Add16~9 ;
wire \Add16~11 ;
wire \Add16~13 ;
wire \Add16~14_combout ;
wire \sig_req_rsc_shift~66_combout ;
wire \Add17~1_combout ;
wire \trk_block:sig_req_rsc_shift[5]~2_combout ;
wire \sig_req_rsc_shift~60_combout ;
wire \sig_req_rsc_shift~67_combout ;
wire \trk_block:sig_req_rsc_shift[7]~q ;
wire \Add18~1 ;
wire \Add18~3 ;
wire \Add18~5 ;
wire \Add18~6_combout ;
wire \trk_block:sig_req_rsc_shift[3]~0_combout ;
wire \Add18~4_combout ;
wire \trk_block:sig_req_rsc_shift[2]~0_combout ;
wire \Add18~2_combout ;
wire \trk_block:sig_req_rsc_shift[1]~0_combout ;
wire \sig_req_rsc_shift~54_combout ;
wire \Add18~0_combout ;
wire \Add16~0_combout ;
wire \sig_req_rsc_shift~55_combout ;
wire \sig_req_rsc_shift~56_combout ;
wire \trk_block:sig_req_rsc_shift[5]~1_combout ;
wire \trk_block:sig_req_rsc_shift[5]~3_combout ;
wire \sig_req_rsc_shift~57_combout ;
wire \trk_block:sig_req_rsc_shift[0]~q ;
wire \Add15~1 ;
wire \Add15~2_combout ;
wire \trk_block:sig_req_rsc_shift[5]~4_combout ;
wire \trk_block:sig_req_rsc_shift[1]~q ;
wire \Add15~3 ;
wire \Add15~4_combout ;
wire \trk_block:sig_req_rsc_shift[2]~q ;
wire \Add15~5 ;
wire \Add15~6_combout ;
wire \trk_block:sig_req_rsc_shift[3]~q ;
wire \LessThan10~1_combout ;
wire \sig_trk_state~106_combout ;
wire \sig_phs_shft_start~0_combout ;
wire \sig_phs_shft_start~q ;
wire \Selector126~0_combout ;
wire \sig_trk_pll_start_reconfig~q ;
wire \seq_pll_start_reconfig~2_combout ;
wire \sig_dgrb_last_state.s_release_admin~q ;
wire \ac_handshake_proc~1_combout ;
wire \seq_pll_select~6_combout ;
wire \seq_pll_select~7_combout ;
wire \v_cdvw_state~457_combout ;
wire \sig_cdvw_state.largest_window_size[5]~q ;
wire \dgrb_ctrl~8_combout ;
wire \v_cdvw_state~458_combout ;
wire \sig_cdvw_state.largest_window_size[4]~q ;
wire \dgrb_ctrl~9_combout ;
wire \v_cdvw_state~459_combout ;
wire \sig_cdvw_state.largest_window_size[3]~q ;
wire \dgrb_ctrl~10_combout ;
wire \v_cdvw_state~460_combout ;
wire \sig_cdvw_state.largest_window_size[2]~q ;
wire \dgrb_ctrl~11_combout ;
wire \dgrb_ctrl~12_combout ;
wire \dgrb_ctrl~13_combout ;
wire \sig_mmc_start~5_combout ;
wire \trk_block:sig_mmc_start~q ;
wire \trk_block:mimic_sample_req:v_echo~q ;
wire \seq_mmc_start~1_combout ;


dffeas \ac_block:sig_doing_rd_count (
	.clk(clk),
	.d(\sig_doing_rd_count~10_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.sload(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.ena(vcc),
	.q(\ac_block:sig_doing_rd_count~q ),
	.prn(vcc));
defparam \ac_block:sig_doing_rd_count .is_wysiwyg = "true";
defparam \ac_block:sig_doing_rd_count .power_up = "low";

cycloneiii_lcell_comb \Add23~0 (
	.dataa(\ac_block:sig_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add23~0_combout ),
	.cout(\Add23~1 ));
defparam \Add23~0 .lut_mask = 16'h55AA;
defparam \Add23~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add23~2 (
	.dataa(\ac_block:sig_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~1 ),
	.combout(\Add23~2_combout ),
	.cout(\Add23~3 ));
defparam \Add23~2 .lut_mask = 16'h5A5F;
defparam \Add23~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add23~4 (
	.dataa(\ac_block:sig_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~3 ),
	.combout(\Add23~4_combout ),
	.cout(\Add23~5 ));
defparam \Add23~4 .lut_mask = 16'h5AAF;
defparam \Add23~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add23~12 (
	.dataa(\ac_block:sig_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~11 ),
	.combout(\Add23~12_combout ),
	.cout(\Add23~13 ));
defparam \Add23~12 .lut_mask = 16'h5AAF;
defparam \Add23~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add23~14 (
	.dataa(\ac_block:sig_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add23~13 ),
	.combout(\Add23~14_combout ),
	.cout());
defparam \Add23~14 .lut_mask = 16'h5A5A;
defparam \Add23~14 .sum_lutc_input = "cin";

dffeas sig_trk_ack(
	.clk(clk),
	.d(\Selector127~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_ack~q ),
	.prn(vcc));
defparam sig_trk_ack.is_wysiwyg = "true";
defparam sig_trk_ack.power_up = "low";

dffeas \trk_block:sig_req_rsc_shift[5] (
	.clk(clk),
	.d(\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.asdata(\Add15~10_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sload(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.ena(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.q(\trk_block:sig_req_rsc_shift[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[5] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[5] .power_up = "low";

dffeas \trk_block:sig_req_rsc_shift[4] (
	.clk(clk),
	.d(\trk_block:sig_req_rsc_shift[4]~0_combout ),
	.asdata(\Add15~8_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sload(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.ena(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.q(\trk_block:sig_req_rsc_shift[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[4] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[4] .power_up = "low";

dffeas \trk_block:sig_mimic_delta[0] (
	.clk(clk),
	.d(\Add11~28_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[0] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[0] .power_up = "low";

cycloneiii_lcell_comb \Add15~0 (
	.dataa(\trk_block:sig_mimic_delta[0]~q ),
	.datab(\trk_block:sig_req_rsc_shift[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add15~0_combout ),
	.cout(\Add15~1 ));
defparam \Add15~0 .lut_mask = 16'h66BB;
defparam \Add15~0 .sum_lutc_input = "datac";

dffeas \trk_block:sig_large_drift_seen (
	.clk(clk),
	.d(\LessThan7~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.ena(vcc),
	.q(\trk_block:sig_large_drift_seen~q ),
	.prn(vcc));
defparam \trk_block:sig_large_drift_seen .is_wysiwyg = "true";
defparam \trk_block:sig_large_drift_seen .power_up = "low";

dffeas \trk_block:sig_mimic_delta[5] (
	.clk(clk),
	.d(\Add11~29_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[5] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[5] .power_up = "low";

dffeas \trk_block:sig_mimic_delta[4] (
	.clk(clk),
	.d(\Add11~30_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[4] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[4] .power_up = "low";

dffeas \trk_block:sig_mimic_delta[3] (
	.clk(clk),
	.d(\Add11~31_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[3] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[3] .power_up = "low";

dffeas \trk_block:sig_mimic_delta[2] (
	.clk(clk),
	.d(\Add11~32_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[2] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[2] .power_up = "low";

dffeas \trk_block:sig_mimic_delta[1] (
	.clk(clk),
	.d(\Add11~33_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[1] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[1] .power_up = "low";

cycloneiii_lcell_comb \Add15~6 (
	.dataa(\trk_block:sig_mimic_delta[3]~q ),
	.datab(\trk_block:sig_req_rsc_shift[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~5 ),
	.combout(\Add15~6_combout ),
	.cout(\Add15~7 ));
defparam \Add15~6 .lut_mask = 16'h967F;
defparam \Add15~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add15~8 (
	.dataa(\trk_block:sig_mimic_delta[4]~q ),
	.datab(\trk_block:sig_req_rsc_shift[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~7 ),
	.combout(\Add15~8_combout ),
	.cout(\Add15~9 ));
defparam \Add15~8 .lut_mask = 16'h96EF;
defparam \Add15~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add15~10 (
	.dataa(\trk_block:sig_mimic_delta[5]~q ),
	.datab(\trk_block:sig_req_rsc_shift[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~9 ),
	.combout(\Add15~10_combout ),
	.cout(\Add15~11 ));
defparam \Add15~10 .lut_mask = 16'h967F;
defparam \Add15~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add15~12 (
	.dataa(\trk_block:sig_mimic_delta[7]~q ),
	.datab(\trk_block:sig_req_rsc_shift[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~11 ),
	.combout(\Add15~12_combout ),
	.cout(\Add15~13 ));
defparam \Add15~12 .lut_mask = 16'h96DF;
defparam \Add15~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~2 (
	.dataa(\trk_block:sig_req_rsc_shift[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~1 ),
	.combout(\Add16~2_combout ),
	.cout(\Add16~3 ));
defparam \Add16~2 .lut_mask = 16'h5A5F;
defparam \Add16~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~4 (
	.dataa(\trk_block:sig_req_rsc_shift[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~3 ),
	.combout(\Add16~4_combout ),
	.cout(\Add16~5 ));
defparam \Add16~4 .lut_mask = 16'h5AAF;
defparam \Add16~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~6 (
	.dataa(\trk_block:sig_req_rsc_shift[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~5 ),
	.combout(\Add16~6_combout ),
	.cout(\Add16~7 ));
defparam \Add16~6 .lut_mask = 16'h5A5F;
defparam \Add16~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~8 (
	.dataa(\trk_block:sig_req_rsc_shift[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~7 ),
	.combout(\Add16~8_combout ),
	.cout(\Add16~9 ));
defparam \Add16~8 .lut_mask = 16'h5AAF;
defparam \Add16~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~10 (
	.dataa(\trk_block:sig_req_rsc_shift[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~9 ),
	.combout(\Add16~10_combout ),
	.cout(\Add16~11 ));
defparam \Add16~10 .lut_mask = 16'h5A5F;
defparam \Add16~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add16~12 (
	.dataa(\trk_block:sig_req_rsc_shift[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add16~11 ),
	.combout(\Add16~12_combout ),
	.cout(\Add16~13 ));
defparam \Add16~12 .lut_mask = 16'h5AAF;
defparam \Add16~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~6 (
	.dataa(\trk_block:sig_req_rsc_shift[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~5 ),
	.combout(\Add18~6_combout ),
	.cout(\Add18~7 ));
defparam \Add18~6 .lut_mask = 16'h5A5F;
defparam \Add18~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~8 (
	.dataa(\trk_block:sig_req_rsc_shift[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~7 ),
	.combout(\Add18~8_combout ),
	.cout(\Add18~9 ));
defparam \Add18~8 .lut_mask = 16'h5AAF;
defparam \Add18~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~10 (
	.dataa(\trk_block:sig_req_rsc_shift[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~9 ),
	.combout(\Add18~10_combout ),
	.cout(\Add18~11 ));
defparam \Add18~10 .lut_mask = 16'h5A5F;
defparam \Add18~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~12 (
	.dataa(\trk_block:sig_req_rsc_shift[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~11 ),
	.combout(\Add18~12_combout ),
	.cout(\Add18~13 ));
defparam \Add18~12 .lut_mask = 16'h5AAF;
defparam \Add18~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[5]~0 (
	.dataa(\Add16~10_combout ),
	.datab(\Add18~10_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[5]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_req_rsc_shift[5]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[4]~0 (
	.dataa(\Add16~8_combout ),
	.datab(\Add18~8_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[4]~0_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[4]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_req_rsc_shift[4]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add15~14 (
	.dataa(\trk_block:sig_mimic_delta[7]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add15~13 ),
	.combout(\Add15~14_combout ),
	.cout());
defparam \Add15~14 .lut_mask = 16'h9696;
defparam \Add15~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~14 (
	.dataa(\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add18~13 ),
	.combout(\Add18~14_combout ),
	.cout());
defparam \Add18~14 .lut_mask = 16'h5A5A;
defparam \Add18~14 .sum_lutc_input = "cin";

dffeas \trk_block:trk_proc:v_remaining_samples[3] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[3]~0_combout ),
	.asdata(\Selector122~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[3]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[3] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[3] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[6] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[6]~0_combout ),
	.asdata(\sig_rsc_drift~40_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[6] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[6] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[5] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[5]~0_combout ),
	.asdata(\sig_rsc_drift~41_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[5] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[5] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[4] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[4]~0_combout ),
	.asdata(\sig_rsc_drift~42_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[4] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[4] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[3] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[3]~0_combout ),
	.asdata(\sig_rsc_drift~43_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[3] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[3] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[2] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[2]~0_combout ),
	.asdata(\sig_rsc_drift~44_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[2] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[2] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[1] (
	.clk(clk),
	.d(\trk_block:sig_rsc_drift[1]~0_combout ),
	.asdata(\sig_rsc_drift~45_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\sig_dgrb_state.s_track~q ),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[1] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[1] .power_up = "low";

cycloneiii_lcell_comb \Add9~0 (
	.dataa(\trk_block:sig_rsc_drift[0]~q ),
	.datab(\cal_codvw_phase[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add9~0_combout ),
	.cout(\Add9~1 ));
defparam \Add9~0 .lut_mask = 16'h66DD;
defparam \Add9~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add9~2 (
	.dataa(\trk_block:sig_rsc_drift[1]~q ),
	.datab(\cal_codvw_phase[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~1 ),
	.combout(\Add9~2_combout ),
	.cout(\Add9~3 ));
defparam \Add9~2 .lut_mask = 16'h967F;
defparam \Add9~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~4 (
	.dataa(\trk_block:sig_rsc_drift[2]~q ),
	.datab(\cal_codvw_phase[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~3 ),
	.combout(\Add9~4_combout ),
	.cout(\Add9~5 ));
defparam \Add9~4 .lut_mask = 16'h96EF;
defparam \Add9~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~6 (
	.dataa(\trk_block:sig_rsc_drift[3]~q ),
	.datab(\cal_codvw_phase[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~5 ),
	.combout(\Add9~6_combout ),
	.cout(\Add9~7 ));
defparam \Add9~6 .lut_mask = 16'h967F;
defparam \Add9~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~8 (
	.dataa(\trk_block:sig_rsc_drift[4]~q ),
	.datab(\cal_codvw_phase[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~7 ),
	.combout(\Add9~8_combout ),
	.cout(\Add9~9 ));
defparam \Add9~8 .lut_mask = 16'h96EF;
defparam \Add9~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~10 (
	.dataa(\trk_block:sig_rsc_drift[5]~q ),
	.datab(\cal_codvw_phase[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~9 ),
	.combout(\Add9~10_combout ),
	.cout(\Add9~11 ));
defparam \Add9~10 .lut_mask = 16'h967F;
defparam \Add9~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~13 (
	.dataa(\trk_block:sig_rsc_drift[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~11 ),
	.combout(),
	.cout(\Add9~13_cout ));
defparam \Add9~13 .lut_mask = 16'h00AF;
defparam \Add9~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~15 (
	.dataa(\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add9~13_cout ),
	.combout(),
	.cout(\Add9~15_cout ));
defparam \Add9~15 .lut_mask = 16'h00AF;
defparam \Add9~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add9~16 (
	.dataa(\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add9~15_cout ),
	.combout(\Add9~16_combout ),
	.cout());
defparam \Add9~16 .lut_mask = 16'h5A5A;
defparam \Add9~16 .sum_lutc_input = "cin";

dffeas \rsc_block:sig_test_dq_expired (
	.clk(clk),
	.d(\sig_test_dq_expired~6_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\rsc_block:sig_test_dq_expired~q ),
	.prn(vcc));
defparam \rsc_block:sig_test_dq_expired .is_wysiwyg = "true";
defparam \rsc_block:sig_test_dq_expired .power_up = "low";

cycloneiii_lcell_comb \Add5~17 (
	.dataa(\Add5~4_combout ),
	.datab(\Add5~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~16 ),
	.combout(\Add5~17_combout ),
	.cout(\Add5~18 ));
defparam \Add5~17 .lut_mask = 16'h96BF;
defparam \Add5~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add5~19 (
	.dataa(\Add5~2_combout ),
	.datab(\Add5~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add5~18 ),
	.combout(\Add5~19_combout ),
	.cout());
defparam \Add5~19 .lut_mask = 16'h9696;
defparam \Add5~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~0 (
	.dataa(\rsc_block:sig_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add6~0_combout ),
	.cout(\Add6~1 ));
defparam \Add6~0 .lut_mask = 16'h55AA;
defparam \Add6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add6~2 (
	.dataa(\rsc_block:sig_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~1 ),
	.combout(\Add6~2_combout ),
	.cout(\Add6~3 ));
defparam \Add6~2 .lut_mask = 16'h5A5F;
defparam \Add6~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~4 (
	.dataa(\rsc_block:sig_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~3 ),
	.combout(\Add6~4_combout ),
	.cout(\Add6~5 ));
defparam \Add6~4 .lut_mask = 16'h5AAF;
defparam \Add6~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~6 (
	.dataa(\rsc_block:sig_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~5 ),
	.combout(\Add6~6_combout ),
	.cout(\Add6~7 ));
defparam \Add6~6 .lut_mask = 16'h5A5F;
defparam \Add6~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~8 (
	.dataa(\rsc_block:sig_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~7 ),
	.combout(\Add6~8_combout ),
	.cout(\Add6~9 ));
defparam \Add6~8 .lut_mask = 16'h5AAF;
defparam \Add6~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~10 (
	.dataa(\rsc_block:sig_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~9 ),
	.combout(\Add6~10_combout ),
	.cout(\Add6~11 ));
defparam \Add6~10 .lut_mask = 16'h5A5F;
defparam \Add6~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~12 (
	.dataa(\rsc_block:sig_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add6~11 ),
	.combout(\Add6~12_combout ),
	.cout(\Add6~13 ));
defparam \Add6~12 .lut_mask = 16'h5AAF;
defparam \Add6~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add6~14 (
	.dataa(\rsc_block:sig_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add6~13 ),
	.combout(\Add6~14_combout ),
	.cout());
defparam \Add6~14 .lut_mask = 16'h5A5A;
defparam \Add6~14 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_bit[0] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[0]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[0] .power_up = "low";

cycloneiii_lcell_comb \Add11~12 (
	.dataa(\trk_block:sig_mimic_cdv[0]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add11~12_combout ),
	.cout(\Add11~13 ));
defparam \Add11~12 .lut_mask = 16'h66BB;
defparam \Add11~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add12~0 (
	.dataa(\trk_block:sig_mimic_delta[7]~q ),
	.datab(\trk_proc~6_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add12~0_combout ),
	.cout(\Add12~1 ));
defparam \Add12~0 .lut_mask = 16'h6677;
defparam \Add12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add12~2 (
	.dataa(\trk_block:sig_mimic_delta[1]~q ),
	.datab(\trk_block:sig_mimic_delta[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add12~1 ),
	.combout(\Add12~2_combout ),
	.cout(\Add12~3 ));
defparam \Add12~2 .lut_mask = 16'h966F;
defparam \Add12~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add12~4 (
	.dataa(\trk_block:sig_mimic_delta[2]~q ),
	.datab(\trk_block:sig_mimic_delta[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add12~3 ),
	.combout(\Add12~4_combout ),
	.cout(\Add12~5 ));
defparam \Add12~4 .lut_mask = 16'h966F;
defparam \Add12~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add12~6 (
	.dataa(\trk_block:sig_mimic_delta[3]~q ),
	.datab(\trk_block:sig_mimic_delta[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add12~5 ),
	.combout(\Add12~6_combout ),
	.cout(\Add12~7 ));
defparam \Add12~6 .lut_mask = 16'h966F;
defparam \Add12~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add12~8 (
	.dataa(\trk_block:sig_mimic_delta[4]~q ),
	.datab(\trk_block:sig_mimic_delta[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add12~7 ),
	.combout(\Add12~8_combout ),
	.cout(\Add12~9 ));
defparam \Add12~8 .lut_mask = 16'h966F;
defparam \Add12~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add12~10 (
	.dataa(\trk_block:sig_mimic_delta[5]~q ),
	.datab(\trk_block:sig_mimic_delta[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add12~9 ),
	.combout(\Add12~10_combout ),
	.cout(\Add12~11 ));
defparam \Add12~10 .lut_mask = 16'h966F;
defparam \Add12~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add12~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add12~11 ),
	.combout(\Add12~12_combout ),
	.cout());
defparam \Add12~12 .lut_mask = 16'h0F0F;
defparam \Add12~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~15 (
	.dataa(\trk_block:sig_mimic_cdv[1]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add11~13 ),
	.combout(\Add11~15_combout ),
	.cout(\Add11~16 ));
defparam \Add11~15 .lut_mask = 16'h96DF;
defparam \Add11~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~17 (
	.dataa(\trk_block:sig_mimic_cdv[2]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add11~16 ),
	.combout(\Add11~17_combout ),
	.cout(\Add11~18 ));
defparam \Add11~17 .lut_mask = 16'h96BF;
defparam \Add11~17 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~19 (
	.dataa(\trk_block:sig_mimic_cdv[3]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add11~18 ),
	.combout(\Add11~19_combout ),
	.cout(\Add11~20 ));
defparam \Add11~19 .lut_mask = 16'h96DF;
defparam \Add11~19 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~21 (
	.dataa(\trk_block:sig_mimic_cdv[4]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add11~20 ),
	.combout(\Add11~21_combout ),
	.cout(\Add11~22 ));
defparam \Add11~21 .lut_mask = 16'h96BF;
defparam \Add11~21 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~23 (
	.dataa(\trk_block:sig_mimic_cdv[5]~q ),
	.datab(\sig_cdvw_state.largest_window_centre[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add11~22 ),
	.combout(\Add11~23_combout ),
	.cout(\Add11~24 ));
defparam \Add11~23 .lut_mask = 16'h96DF;
defparam \Add11~23 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add11~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add11~24 ),
	.combout(\Add11~25_combout ),
	.cout());
defparam \Add11~25 .lut_mask = 16'hF0F0;
defparam \Add11~25 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add10~0_combout ),
	.cout(\Add10~1 ));
defparam \Add10~0 .lut_mask = 16'h55AA;
defparam \Add10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add10~2 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~1 ),
	.combout(\Add10~2_combout ),
	.cout(\Add10~3 ));
defparam \Add10~2 .lut_mask = 16'h5A5F;
defparam \Add10~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~4 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~3 ),
	.combout(\Add10~4_combout ),
	.cout(\Add10~5 ));
defparam \Add10~4 .lut_mask = 16'h5AAF;
defparam \Add10~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~6 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~5 ),
	.combout(\Add10~6_combout ),
	.cout(\Add10~7 ));
defparam \Add10~6 .lut_mask = 16'h5A5F;
defparam \Add10~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~8 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~7 ),
	.combout(\Add10~8_combout ),
	.cout(\Add10~9 ));
defparam \Add10~8 .lut_mask = 16'h5AAF;
defparam \Add10~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~10 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~9 ),
	.combout(\Add10~10_combout ),
	.cout(\Add10~11 ));
defparam \Add10~10 .lut_mask = 16'h5A5F;
defparam \Add10~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~12 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~11 ),
	.combout(\Add10~12_combout ),
	.cout(\Add10~13 ));
defparam \Add10~12 .lut_mask = 16'h5AAF;
defparam \Add10~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add10~14 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add10~13 ),
	.combout(\Add10~14_combout ),
	.cout());
defparam \Add10~14 .lut_mask = 16'h5A5A;
defparam \Add10~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[3]~0 (
	.dataa(\Add10~6_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[3]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[3]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[3]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~3 (
	.dataa(\trk_block:sig_rsc_drift[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add17~3_cout ));
defparam \Add17~3 .lut_mask = 16'h0055;
defparam \Add17~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~4 (
	.dataa(\trk_block:sig_rsc_drift[1]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~3_cout ),
	.combout(\Add17~4_combout ),
	.cout(\Add17~5 ));
defparam \Add17~4 .lut_mask = 16'h967F;
defparam \Add17~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~6 (
	.dataa(\trk_block:sig_rsc_drift[2]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~5 ),
	.combout(\Add17~6_combout ),
	.cout(\Add17~7 ));
defparam \Add17~6 .lut_mask = 16'h96EF;
defparam \Add17~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~8 (
	.dataa(\trk_block:sig_rsc_drift[3]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~7 ),
	.combout(\Add17~8_combout ),
	.cout(\Add17~9 ));
defparam \Add17~8 .lut_mask = 16'h967F;
defparam \Add17~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~10 (
	.dataa(\trk_block:sig_rsc_drift[4]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~9 ),
	.combout(\Add17~10_combout ),
	.cout(\Add17~11 ));
defparam \Add17~10 .lut_mask = 16'h96EF;
defparam \Add17~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~12 (
	.dataa(\trk_block:sig_rsc_drift[5]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~11 ),
	.combout(\Add17~12_combout ),
	.cout(\Add17~13 ));
defparam \Add17~12 .lut_mask = 16'h967F;
defparam \Add17~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~14 (
	.dataa(\trk_block:sig_rsc_drift[6]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add17~13 ),
	.combout(\Add17~14_combout ),
	.cout(\Add17~15 ));
defparam \Add17~14 .lut_mask = 16'h96EF;
defparam \Add17~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add17~16 (
	.dataa(\trk_block:sig_rsc_drift[7]~q ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add17~15 ),
	.combout(\Add17~16_combout ),
	.cout());
defparam \Add17~16 .lut_mask = 16'h9696;
defparam \Add17~16 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[6]~0 (
	.dataa(\Selector95~0_combout ),
	.datab(\Add17~21_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[6]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[6]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[6]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[5]~0 (
	.dataa(\Selector96~0_combout ),
	.datab(\Add17~22_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[5]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[5]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[5]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[4]~0 (
	.dataa(\Selector97~0_combout ),
	.datab(\Add17~23_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[4]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[4]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[4]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[3]~0 (
	.dataa(\Selector98~0_combout ),
	.datab(\Add17~24_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[3]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[3]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[2]~0 (
	.dataa(\Selector99~0_combout ),
	.datab(\Add17~25_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[2]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[2]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_rsc_drift[1]~0 (
	.dataa(\Selector100~0_combout ),
	.datab(\Add17~26_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\trk_block:sig_rsc_drift[1]~0_combout ),
	.cout());
defparam \trk_block:sig_rsc_drift[1]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_rsc_drift[1]~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.current_window_centre[5] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[5]~16_combout ),
	.asdata(\sig_cdvw_state.current_bit[5]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[5] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[4] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[4]~14_combout ),
	.asdata(\sig_cdvw_state.current_bit[4]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[4] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[3] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[3]~12_combout ),
	.asdata(\sig_cdvw_state.current_bit[3]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[3] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[2] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[2]~10_combout ),
	.asdata(\sig_cdvw_state.current_bit[2]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[2] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[1] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[1]~8_combout ),
	.asdata(\sig_cdvw_state.current_bit[1]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[1] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[0] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[0]~6_combout ),
	.asdata(\sig_cdvw_state.current_bit[0]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.sload(\find_centre_of_largest_data_valid_window~6_combout ),
	.ena(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.q(\sig_cdvw_state.current_window_centre[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[0] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[0]~6 (
	.dataa(\sig_cdvw_state.current_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_bit[0]~6_combout ),
	.cout(\sig_cdvw_state.current_bit[0]~7 ));
defparam \sig_cdvw_state.current_bit[0]~6 .lut_mask = 16'h55AA;
defparam \sig_cdvw_state.current_bit[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[0]~6 (
	.dataa(\sig_cdvw_state.current_window_centre[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[0]~6_combout ),
	.cout(\sig_cdvw_state.current_window_centre[0]~7 ));
defparam \sig_cdvw_state.current_window_centre[0]~6 .lut_mask = 16'h55AA;
defparam \sig_cdvw_state.current_window_centre[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[1]~8 (
	.dataa(\sig_cdvw_state.current_window_centre[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_centre[0]~7 ),
	.combout(\sig_cdvw_state.current_window_centre[1]~8_combout ),
	.cout(\sig_cdvw_state.current_window_centre[1]~9 ));
defparam \sig_cdvw_state.current_window_centre[1]~8 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_window_centre[1]~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[2]~10 (
	.dataa(\sig_cdvw_state.current_window_centre[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_centre[1]~9 ),
	.combout(\sig_cdvw_state.current_window_centre[2]~10_combout ),
	.cout(\sig_cdvw_state.current_window_centre[2]~11 ));
defparam \sig_cdvw_state.current_window_centre[2]~10 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_window_centre[2]~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[3]~12 (
	.dataa(\sig_cdvw_state.current_window_centre[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_centre[2]~11 ),
	.combout(\sig_cdvw_state.current_window_centre[3]~12_combout ),
	.cout(\sig_cdvw_state.current_window_centre[3]~13 ));
defparam \sig_cdvw_state.current_window_centre[3]~12 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_window_centre[3]~12 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[4]~14 (
	.dataa(\sig_cdvw_state.current_window_centre[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_centre[3]~13 ),
	.combout(\sig_cdvw_state.current_window_centre[4]~14_combout ),
	.cout(\sig_cdvw_state.current_window_centre[4]~15 ));
defparam \sig_cdvw_state.current_window_centre[4]~14 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_window_centre[4]~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~16 (
	.dataa(\sig_cdvw_state.current_window_centre[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sig_cdvw_state.current_window_centre[4]~15 ),
	.combout(\sig_cdvw_state.current_window_centre[5]~16_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~16 .lut_mask = 16'h5A5A;
defparam \sig_cdvw_state.current_window_centre[5]~16 .sum_lutc_input = "cin";

dffeas sig_rsc_cdvw_phase(
	.clk(clk),
	.d(\sig_rsc_cdvw_phase~5_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\sig_rsc_cdvw_phase~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_phase.is_wysiwyg = "true";
defparam sig_rsc_cdvw_phase.power_up = "low";

dffeas \ac_block:sig_count[7] (
	.clk(clk),
	.d(\Selector166~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~7_combout ),
	.q(\ac_block:sig_count[7]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[7] .is_wysiwyg = "true";
defparam \ac_block:sig_count[7] .power_up = "low";

cycloneiii_lcell_comb \Selector140~6 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\Selector140~6_combout ),
	.cout());
defparam \Selector140~6 .lut_mask = 16'hEEFF;
defparam \Selector140~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[12]~0 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(\Equal13~1_combout ),
	.datad(\Selector174~0_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~0_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[12]~0 .lut_mask = 16'h8BFF;
defparam \sig_addr_cmd[0].addr[12]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[12]~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~1_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[12]~1 .lut_mask = 16'hEFFF;
defparam \sig_addr_cmd[0].addr[12]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[7]~3 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datab(\Equal13~1_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~3_combout ),
	.cout());
defparam \ac_block:sig_count[7]~3 .lut_mask = 16'hEEFF;
defparam \ac_block:sig_count[7]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector166~0 (
	.dataa(\ac_block:sig_count[7]~2_combout ),
	.datab(\Add23~14_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_count[7]~5_combout ),
	.cin(gnd),
	.combout(\Selector166~0_combout ),
	.cout());
defparam \Selector166~0 .lut_mask = 16'hEEFF;
defparam \Selector166~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[7]~6 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(dgb_ac_access_gnt_r),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~6_combout ),
	.cout());
defparam \ac_block:sig_count[7]~6 .lut_mask = 16'hEFFF;
defparam \ac_block:sig_count[7]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector170~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\Selector170~0_combout ),
	.cout());
defparam \Selector170~0 .lut_mask = 16'hEFFF;
defparam \Selector170~0 .sum_lutc_input = "datac";

dffeas \sig_ac_req.s_ac_read_wd_lat (
	.clk(clk),
	.d(\Selector26~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_wd_lat .power_up = "low";

cycloneiii_lcell_comb \WideOr26~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datad(\sig_ac_req.s_ac_read_wd_lat~q ),
	.cin(gnd),
	.combout(\WideOr26~0_combout ),
	.cout());
defparam \WideOr26~0 .lut_mask = 16'h6996;
defparam \WideOr26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[5]~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\Equal13~1_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[5]~1_combout ),
	.cout());
defparam \ac_block:sig_count[5]~1 .lut_mask = 16'hEEFF;
defparam \ac_block:sig_count[5]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~2 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\Selector169~1_combout ),
	.datac(\sig_count~171_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\Selector169~2_combout ),
	.cout());
defparam \Selector169~2 .lut_mask = 16'hEFFF;
defparam \Selector169~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~3 (
	.dataa(\Selector169~2_combout ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(\Selector174~2_combout ),
	.cin(gnd),
	.combout(\Selector169~3_combout ),
	.cout());
defparam \Selector169~3 .lut_mask = 16'hFFFE;
defparam \Selector169~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~4 (
	.dataa(\ac_block:sig_count[7]~0_combout ),
	.datab(\ac_block:sig_count[7]~1_combout ),
	.datac(\ac_block:sig_count[4]~q ),
	.datad(\Selector169~3_combout ),
	.cin(gnd),
	.combout(\Selector169~4_combout ),
	.cout());
defparam \Selector169~4 .lut_mask = 16'hFFFE;
defparam \Selector169~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_doing_rd_count~10 (
	.dataa(\Equal13~0_combout ),
	.datab(\sig_count~171_combout ),
	.datac(\ac_block:sig_count[0]~q ),
	.datad(\ac_block:sig_count[1]~q ),
	.cin(gnd),
	.combout(\sig_doing_rd_count~10_combout ),
	.cout());
defparam \sig_doing_rd_count~10 .lut_mask = 16'hEFFF;
defparam \sig_doing_rd_count~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector25~0 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_state.s_wait_admin~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
defparam \Selector25~0 .lut_mask = 16'hFEFE;
defparam \Selector25~0 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_poa_cal (
	.clk(clk),
	.d(\sig_dgrb_state~275_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_poa_cal~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_poa_cal .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_poa_cal .power_up = "low";

cycloneiii_lcell_comb \Selector26~0 (
	.dataa(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(\sig_ac_req.s_ac_read_wd_lat~q ),
	.datac(\Selector25~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hFEFE;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector21~0 (
	.dataa(\Selector25~1_combout ),
	.datab(\Selector23~0_combout ),
	.datac(\sig_ac_req.s_ac_idle~q ),
	.datad(\sig_rsc_ac_access_req~q ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
defparam \Selector21~0 .lut_mask = 16'hEFFF;
defparam \Selector21~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~244 (
	.dataa(\sig_dgrb_state.s_idle~q ),
	.datab(\sig_dgrb_state~242_combout ),
	.datac(\sig_dgrb_state~243_combout ),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\sig_dgrb_state~244_combout ),
	.cout());
defparam \sig_dgrb_state~244 .lut_mask = 16'hD8FF;
defparam \sig_dgrb_state~244 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~245 (
	.dataa(rdata_valid[0]),
	.datab(\sig_dgrb_state.s_adv_rd_lat~q ),
	.datac(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~245_combout ),
	.cout());
defparam \sig_dgrb_state~245 .lut_mask = 16'hFEFF;
defparam \sig_dgrb_state~245 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~248 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datac(\sig_dgrb_state.s_poa_cal~q ),
	.datad(\sig_dgrb_state.s_adv_rd_lat~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~248_combout ),
	.cout());
defparam \sig_dgrb_state~248 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~248 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~249 (
	.dataa(\sig_dgrb_state.s_idle~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~249_combout ),
	.cout());
defparam \sig_dgrb_state~249 .lut_mask = 16'hAAFF;
defparam \sig_dgrb_state~249 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~250 (
	.dataa(\sig_dgrb_state~244_combout ),
	.datab(\sig_dgrb_state~247_combout ),
	.datac(\sig_dgrb_state~248_combout ),
	.datad(\sig_dgrb_state~249_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~250_combout ),
	.cout());
defparam \sig_dgrb_state~250 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~250 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~252 (
	.dataa(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datab(\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~252_combout ),
	.cout());
defparam \sig_dgrb_state~252 .lut_mask = 16'hEEEE;
defparam \sig_dgrb_state~252 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~253 (
	.dataa(\sig_dgrb_state~251_combout ),
	.datab(\sig_dgrb_state~252_combout ),
	.datac(ac_muxctrl_broadcast_rcommand_req),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~253_combout ),
	.cout());
defparam \sig_dgrb_state~253 .lut_mask = 16'hFAFC;
defparam \sig_dgrb_state~253 .sum_lutc_input = "datac";

dffeas \trk_block:sig_req_rsc_shift[6] (
	.clk(clk),
	.d(\sig_req_rsc_shift~62_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_req_rsc_shift[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[6] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[6] .power_up = "low";

cycloneiii_lcell_comb \LessThan10~0 (
	.dataa(\trk_block:sig_req_rsc_shift[0]~q ),
	.datab(\trk_block:sig_req_rsc_shift[6]~q ),
	.datac(\trk_block:sig_req_rsc_shift[5]~q ),
	.datad(\trk_block:sig_req_rsc_shift[4]~q ),
	.cin(gnd),
	.combout(\LessThan10~0_combout ),
	.cout());
defparam \LessThan10~0 .lut_mask = 16'hBFFF;
defparam \LessThan10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan10~2 (
	.dataa(\LessThan10~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\LessThan10~2_combout ),
	.cout());
defparam \LessThan10~2 .lut_mask = 16'hAAFF;
defparam \LessThan10~2 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rewind_direction (
	.clk(clk),
	.d(\sig_rewind_direction~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rewind_direction~q ),
	.prn(vcc));
defparam \rsc_block:sig_rewind_direction .is_wysiwyg = "true";
defparam \rsc_block:sig_rewind_direction .power_up = "low";

dffeas \rsc_block:sig_num_phase_shifts[5] (
	.clk(clk),
	.d(\Add5~21_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[5]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[5] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[5] .power_up = "low";

dffeas \rsc_block:sig_count[7] (
	.clk(clk),
	.d(\Selector39~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[6]~4_combout ),
	.q(\rsc_block:sig_count[7]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[7] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[7] .power_up = "low";

dffeas \rsc_block:sig_count[6] (
	.clk(clk),
	.d(\Selector40~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[6]~4_combout ),
	.q(\rsc_block:sig_count[6]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[6] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[6] .power_up = "low";

dffeas \rsc_block:sig_count[5] (
	.clk(clk),
	.d(\Selector41~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[5]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[5] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[5] .power_up = "low";

dffeas \rsc_block:sig_count[4] (
	.clk(clk),
	.d(\Selector42~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[4]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[4] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[4] .power_up = "low";

cycloneiii_lcell_comb \Equal7~0 (
	.dataa(\rsc_block:sig_count[7]~q ),
	.datab(\rsc_block:sig_count[6]~q ),
	.datac(\rsc_block:sig_count[5]~q ),
	.datad(\rsc_block:sig_count[4]~q ),
	.cin(gnd),
	.combout(\Equal7~0_combout ),
	.cout());
defparam \Equal7~0 .lut_mask = 16'h7FFF;
defparam \Equal7~0 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_count[3] (
	.clk(clk),
	.d(\Selector43~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[3]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[3] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[3] .power_up = "low";

dffeas \rsc_block:sig_count[2] (
	.clk(clk),
	.d(\Selector44~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[2]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[2] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[2] .power_up = "low";

dffeas \rsc_block:sig_count[1] (
	.clk(clk),
	.d(\Selector45~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[1]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[1] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[1] .power_up = "low";

cycloneiii_lcell_comb \Equal7~1 (
	.dataa(\Equal7~0_combout ),
	.datab(\rsc_block:sig_count[3]~q ),
	.datac(\rsc_block:sig_count[2]~q ),
	.datad(\rsc_block:sig_count[1]~q ),
	.cin(gnd),
	.combout(\Equal7~1_combout ),
	.cout());
defparam \Equal7~1 .lut_mask = 16'hBFFF;
defparam \Equal7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector59~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datab(\Selector69~0_combout ),
	.datac(\Equal7~2_combout ),
	.datad(\sig_phs_shft_start~q ),
	.cin(gnd),
	.combout(\Selector59~1_combout ),
	.cout());
defparam \Selector59~1 .lut_mask = 16'hEFFF;
defparam \Selector59~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~266 (
	.dataa(\dgrb_state_proc~4_combout ),
	.datab(\sig_dgrb_state~243_combout ),
	.datac(\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~266_combout ),
	.cout());
defparam \sig_dgrb_state~266 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~266 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_cdvw_wait (
	.clk(clk),
	.d(\Selector56~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_wait .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_wait .power_up = "low";

dffeas \ctrl_dgrb_r.command.cmd_poa (
	.clk(clk),
	.d(Selector52),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_poa~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_poa .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_poa .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~275 (
	.dataa(\sig_dgrb_state.s_wait_admin~q ),
	.datab(\dgrb_state_proc~4_combout ),
	.datac(\ctrl_dgrb_r.command.cmd_poa~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~275_combout ),
	.cout());
defparam \sig_dgrb_state~275 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~275 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~276 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_dgrb_state.s_poa_cal~q ),
	.datac(\sig_poa_ack~q ),
	.datad(\sig_trk_ack~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~276_combout ),
	.cout());
defparam \sig_dgrb_state~276 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~276 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_complete (
	.clk(clk),
	.d(\sig_trk_state~120_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_complete~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_complete .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_complete .power_up = "low";

cycloneiii_lcell_comb \Selector127~0 (
	.dataa(\trk_block:sig_trk_state.s_trk_complete~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\sig_cdvw_state.status.valid_result~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\Selector127~0_combout ),
	.cout());
defparam \Selector127~0 .lut_mask = 16'hEFFF;
defparam \Selector127~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~58 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~58_combout ),
	.cout());
defparam \sig_req_rsc_shift~58 .lut_mask = 16'hFEFE;
defparam \sig_req_rsc_shift~58 .sum_lutc_input = "datac";

dffeas \trk_block:sig_mimic_delta[7] (
	.clk(clk),
	.d(\Add11~27_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Add11~14_combout ),
	.q(\trk_block:sig_mimic_delta[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[7] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[7] .power_up = "low";

cycloneiii_lcell_comb \sig_req_rsc_shift~59 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~59_combout ),
	.cout());
defparam \sig_req_rsc_shift~59 .lut_mask = 16'hEEFF;
defparam \sig_req_rsc_shift~59 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~61 (
	.dataa(\sig_req_rsc_shift~59_combout ),
	.datab(\trk_block:sig_req_rsc_shift[6]~q ),
	.datac(\sig_req_rsc_shift~60_combout ),
	.datad(\sig_req_rsc_shift~68_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~61_combout ),
	.cout());
defparam \sig_req_rsc_shift~61 .lut_mask = 16'hFFFE;
defparam \sig_req_rsc_shift~61 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~62 (
	.dataa(\sig_req_rsc_shift~58_combout ),
	.datab(\trk_block:sig_large_drift_seen~q ),
	.datac(\Add15~12_combout ),
	.datad(\sig_req_rsc_shift~61_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~62_combout ),
	.cout());
defparam \sig_req_rsc_shift~62 .lut_mask = 16'hFFBE;
defparam \sig_req_rsc_shift~62 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~63 (
	.dataa(\trk_block:sig_mimic_delta[7]~q ),
	.datab(\Add15~12_combout ),
	.datac(\Add15~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~63_combout ),
	.cout());
defparam \sig_req_rsc_shift~63 .lut_mask = 16'h9696;
defparam \sig_req_rsc_shift~63 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~64 (
	.dataa(\sig_req_rsc_shift~58_combout ),
	.datab(\sig_req_rsc_shift~63_combout ),
	.datac(\Add15~14_combout ),
	.datad(\trk_block:sig_large_drift_seen~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~64_combout ),
	.cout());
defparam \sig_req_rsc_shift~64 .lut_mask = 16'hFAFC;
defparam \sig_req_rsc_shift~64 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~65 (
	.dataa(\sig_req_rsc_shift~64_combout ),
	.datab(\sig_req_rsc_shift~59_combout ),
	.datac(\Add18~14_combout ),
	.datad(\LessThan10~2_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~65_combout ),
	.cout());
defparam \sig_req_rsc_shift~65 .lut_mask = 16'hFEFF;
defparam \sig_req_rsc_shift~65 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[6] (
	.clk(clk),
	.d(\Selector119~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[6]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[6] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[6] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[7] (
	.clk(clk),
	.d(\Add17~20_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[7] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[7] .power_up = "low";

dffeas \cal_codvw_phase[5] (
	.clk(clk),
	.d(\Selector69~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[5]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[5] .is_wysiwyg = "true";
defparam \cal_codvw_phase[5] .power_up = "low";

dffeas \cal_codvw_phase[4] (
	.clk(clk),
	.d(\Selector70~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[4]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[4] .is_wysiwyg = "true";
defparam \cal_codvw_phase[4] .power_up = "low";

dffeas \cal_codvw_phase[3] (
	.clk(clk),
	.d(\Selector71~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[3]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[3] .is_wysiwyg = "true";
defparam \cal_codvw_phase[3] .power_up = "low";

dffeas \cal_codvw_phase[2] (
	.clk(clk),
	.d(\Selector72~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[2]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[2] .is_wysiwyg = "true";
defparam \cal_codvw_phase[2] .power_up = "low";

dffeas \cal_codvw_phase[1] (
	.clk(clk),
	.d(\Selector73~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[1]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[1] .is_wysiwyg = "true";
defparam \cal_codvw_phase[1] .power_up = "low";

dffeas \trk_block:sig_rsc_drift[0] (
	.clk(clk),
	.d(\Add17~27_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[0] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[0] .power_up = "low";

cycloneiii_lcell_comb \sig_rewind_direction~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datab(\Add9~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rewind_direction~1_combout ),
	.cout());
defparam \sig_rewind_direction~1 .lut_mask = 16'hEEEE;
defparam \sig_rewind_direction~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\Add5~1_combout ),
	.cout());
defparam \Add5~1 .lut_mask = 16'hFEFF;
defparam \Add5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~2 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[5]~q ),
	.datad(\Add9~10_combout ),
	.cin(gnd),
	.combout(\Add5~2_combout ),
	.cout());
defparam \Add5~2 .lut_mask = 16'h8BFF;
defparam \Add5~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~4 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[4]~q ),
	.datad(\Add9~8_combout ),
	.cin(gnd),
	.combout(\Add5~4_combout ),
	.cout());
defparam \Add5~4 .lut_mask = 16'h8BFF;
defparam \Add5~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~5 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[3]~q ),
	.datad(\Add9~6_combout ),
	.cin(gnd),
	.combout(\Add5~5_combout ),
	.cout());
defparam \Add5~5 .lut_mask = 16'h8BFF;
defparam \Add5~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~6 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[2]~q ),
	.datad(\Add9~4_combout ),
	.cin(gnd),
	.combout(\Add5~6_combout ),
	.cout());
defparam \Add5~6 .lut_mask = 16'h8BFF;
defparam \Add5~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~7 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[1]~q ),
	.datad(\Add9~2_combout ),
	.cin(gnd),
	.combout(\Add5~7_combout ),
	.cout());
defparam \Add5~7 .lut_mask = 16'h8BFF;
defparam \Add5~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~21 (
	.dataa(\Add9~10_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~19_combout ),
	.cin(gnd),
	.combout(\Add5~21_combout ),
	.cout());
defparam \Add5~21 .lut_mask = 16'h47FF;
defparam \Add5~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector48~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_phs_shft_end~q ),
	.cin(gnd),
	.combout(\Selector48~0_combout ),
	.cout());
defparam \Selector48~0 .lut_mask = 16'hAAFF;
defparam \Selector48~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector57~0 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_read_mtp~q ),
	.cin(gnd),
	.combout(\Selector57~0_combout ),
	.cout());
defparam \Selector57~0 .lut_mask = 16'hEEFF;
defparam \Selector57~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~0 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datac(gnd),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~0_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~0 .lut_mask = 16'hAACC;
defparam \rsc_block:sig_count[6]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~2 (
	.dataa(\WideOr13~0_combout ),
	.datab(\rsc_block:sig_count[6]~0_combout ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~2_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~2 .lut_mask = 16'hBFFF;
defparam \rsc_block:sig_count[6]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector39~0 (
	.dataa(\Add6~14_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_count[6]~2_combout ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
defparam \Selector39~0 .lut_mask = 16'hAAFF;
defparam \Selector39~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~3 (
	.dataa(\sig_dimm_driving_dq~q ),
	.datab(\rsc_proc~1_combout ),
	.datac(\Equal7~2_combout ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~3_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~3 .lut_mask = 16'hFAFC;
defparam \rsc_block:sig_count[6]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~4 (
	.dataa(\rsc_block:sig_count[6]~3_combout ),
	.datab(\rsc_block:sig_count[6]~0_combout ),
	.datac(\WideOr13~0_combout ),
	.datad(\rsc_block:sig_count[5]~0_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~4_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~4 .lut_mask = 16'hFF7F;
defparam \rsc_block:sig_count[6]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector40~0 (
	.dataa(\Add6~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_count[6]~2_combout ),
	.cin(gnd),
	.combout(\Selector40~0_combout ),
	.cout());
defparam \Selector40~0 .lut_mask = 16'hAAFF;
defparam \Selector40~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[5] (
	.clk(clk),
	.d(\v_cdvw_state~434_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[5] .power_up = "low";

cycloneiii_lcell_comb \Selector41~0 (
	.dataa(\sig_cdvw_state.largest_window_centre[5]~q ),
	.datab(\Add6~10_combout ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\rsc_block:sig_count[5]~2_combout ),
	.cin(gnd),
	.combout(\Selector41~0_combout ),
	.cout());
defparam \Selector41~0 .lut_mask = 16'hACFF;
defparam \Selector41~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~2 (
	.dataa(\rsc_block:sig_count[6]~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(\Add6~8_combout ),
	.datad(\rsc_block:sig_count[5]~1_combout ),
	.cin(gnd),
	.combout(\Selector42~2_combout ),
	.cout());
defparam \Selector42~2 .lut_mask = 16'hFEFF;
defparam \Selector42~2 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[4] (
	.clk(clk),
	.d(\v_cdvw_state~435_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[4] .power_up = "low";

cycloneiii_lcell_comb \Selector43~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(\rsc_block:sig_count[5]~1_combout ),
	.datac(\Add6~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector43~0_combout ),
	.cout());
defparam \Selector43~0 .lut_mask = 16'hFEFE;
defparam \Selector43~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[3] (
	.clk(clk),
	.d(\v_cdvw_state~436_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[3] .power_up = "low";

cycloneiii_lcell_comb \Selector43~1 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.cin(gnd),
	.combout(\Selector43~1_combout ),
	.cout());
defparam \Selector43~1 .lut_mask = 16'hEFFF;
defparam \Selector43~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector43~2 (
	.dataa(\Selector43~0_combout ),
	.datab(\sig_cdvw_state.largest_window_centre[3]~q ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\Selector43~1_combout ),
	.cin(gnd),
	.combout(\Selector43~2_combout ),
	.cout());
defparam \Selector43~2 .lut_mask = 16'hACFF;
defparam \Selector43~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector44~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(\rsc_block:sig_count[5]~1_combout ),
	.datac(\Add6~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector44~0_combout ),
	.cout());
defparam \Selector44~0 .lut_mask = 16'hFEFE;
defparam \Selector44~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[2] (
	.clk(clk),
	.d(\v_cdvw_state~437_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[2] .power_up = "low";

cycloneiii_lcell_comb \Selector44~1 (
	.dataa(\Selector44~0_combout ),
	.datab(\sig_cdvw_state.largest_window_centre[2]~q ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\Selector43~1_combout ),
	.cin(gnd),
	.combout(\Selector44~1_combout ),
	.cout());
defparam \Selector44~1 .lut_mask = 16'hACFF;
defparam \Selector44~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector45~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(\rsc_block:sig_count[5]~1_combout ),
	.datac(\Add6~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector45~0_combout ),
	.cout());
defparam \Selector45~0 .lut_mask = 16'hFEFE;
defparam \Selector45~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[1] (
	.clk(clk),
	.d(\v_cdvw_state~438_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[1] .power_up = "low";

cycloneiii_lcell_comb \Selector45~1 (
	.dataa(\Selector45~0_combout ),
	.datab(\sig_cdvw_state.largest_window_centre[1]~q ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\Selector43~1_combout ),
	.cin(gnd),
	.combout(\Selector45~1_combout ),
	.cout());
defparam \Selector45~1 .lut_mask = 16'hACFF;
defparam \Selector45~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector56~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\Selector56~0_combout ),
	.cout());
defparam \Selector56~0 .lut_mask = 16'hFFFE;
defparam \Selector56~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \find_centre_of_largest_data_valid_window~5 (
	.dataa(\sig_cdvw_state.current_bit[0]~q ),
	.datab(\sig_cdvw_state.current_bit[1]~q ),
	.datac(\sig_cdvw_state.current_bit[2]~q ),
	.datad(\sig_cdvw_state.current_bit[3]~q ),
	.cin(gnd),
	.combout(\find_centre_of_largest_data_valid_window~5_combout ),
	.cout());
defparam \find_centre_of_largest_data_valid_window~5 .lut_mask = 16'h7FFF;
defparam \find_centre_of_largest_data_valid_window~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \find_centre_of_largest_data_valid_window~0 (
	.dataa(\find_centre_of_largest_data_valid_window~5_combout ),
	.datab(\sig_cdvw_state.current_bit[4]~q ),
	.datac(\sig_cdvw_state.current_bit[5]~q ),
	.datad(\sig_cdvw_state.found_a_good_edge~q ),
	.cin(gnd),
	.combout(\find_centre_of_largest_data_valid_window~0_combout ),
	.cout());
defparam \find_centre_of_largest_data_valid_window~0 .lut_mask = 16'hBFFF;
defparam \find_centre_of_largest_data_valid_window~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_good_edge[2] (
	.clk(clk),
	.d(\v_cdvw_state~441_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[2] .power_up = "low";

dffeas \sig_cdvw_state.first_good_edge[5] (
	.clk(clk),
	.d(\v_cdvw_state~442_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[5] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~424 (
	.dataa(\sig_cdvw_state.current_bit[2]~q ),
	.datab(\sig_cdvw_state.first_good_edge[2]~q ),
	.datac(\sig_cdvw_state.current_bit[5]~q ),
	.datad(\sig_cdvw_state.first_good_edge[5]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~424_combout ),
	.cout());
defparam \v_cdvw_state~424 .lut_mask = 16'h6996;
defparam \v_cdvw_state~424 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.invalid_phase_seen (
	.clk(clk),
	.d(\v_cdvw_state~447_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.invalid_phase_seen~q ),
	.prn(vcc));
defparam \sig_cdvw_state.invalid_phase_seen .is_wysiwyg = "true";
defparam \sig_cdvw_state.invalid_phase_seen .power_up = "low";

dffeas \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm (
	.clk(clk),
	.d(\Selector50~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm .power_up = "low";

cycloneiii_lcell_comb \Selector51~2 (
	.dataa(\sig_dimm_driving_dq~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.datac(\Selector51~1_combout ),
	.datad(\rsc_block:sig_chkd_all_dq_pins~q ),
	.cin(gnd),
	.combout(\Selector51~2_combout ),
	.cout());
defparam \Selector51~2 .lut_mask = 16'hFEFF;
defparam \Selector51~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~116 (
	.dataa(\trk_block:sig_trk_state.s_trk_complete~q ),
	.datab(\sig_cdvw_state.status.calculating~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(\trk_block:sig_mimic_cdv_found~q ),
	.cin(gnd),
	.combout(\sig_trk_state~116_combout ),
	.cout());
defparam \sig_trk_state~116 .lut_mask = 16'hBEFF;
defparam \sig_trk_state~116 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~120 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_state~116_combout ),
	.datac(\sig_trk_state~119_combout ),
	.datad(\sig_trk_state~108_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~120_combout ),
	.cout());
defparam \sig_trk_state~120 .lut_mask = 16'hFEFF;
defparam \sig_trk_state~120 .sum_lutc_input = "datac";

dffeas \trk_block:sig_mimic_cdv[0] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[0] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[0] .power_up = "low";

cycloneiii_lcell_comb \Add11~14 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_mimic_cdv[0]~0_combout ),
	.datac(\Selector93~0_combout ),
	.datad(\trk_block:sig_mimic_cdv_found~q ),
	.cin(gnd),
	.combout(\Add11~14_combout ),
	.cout());
defparam \Add11~14 .lut_mask = 16'hEFFF;
defparam \Add11~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_proc~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\trk_block:sig_mimic_delta[7]~q ),
	.datad(\trk_block:sig_mimic_delta[0]~q ),
	.cin(gnd),
	.combout(\trk_proc~6_combout ),
	.cout());
defparam \trk_proc~6 .lut_mask = 16'h0FF0;
defparam \trk_proc~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan7~0 (
	.dataa(\Add12~0_combout ),
	.datab(\Add12~2_combout ),
	.datac(\Add12~4_combout ),
	.datad(\Add12~6_combout ),
	.cin(gnd),
	.combout(\LessThan7~0_combout ),
	.cout());
defparam \LessThan7~0 .lut_mask = 16'hFFFE;
defparam \LessThan7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \LessThan7~1 (
	.dataa(\Add12~12_combout ),
	.datab(\Add12~10_combout ),
	.datac(\Add12~8_combout ),
	.datad(\LessThan7~0_combout ),
	.cin(gnd),
	.combout(\LessThan7~1_combout ),
	.cout());
defparam \LessThan7~1 .lut_mask = 16'hFFFE;
defparam \LessThan7~1 .sum_lutc_input = "datac";

dffeas \trk_block:sig_mimic_cdv[5] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[5] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[5] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[4] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[4] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[4] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[3] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[3] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[3] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[2] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[2] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[2] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[1] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.q(\trk_block:sig_mimic_cdv[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[1] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[1] .power_up = "low";

cycloneiii_lcell_comb \Add11~27 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(\trk_block:sig_mimic_cdv[0]~0_combout ),
	.datad(\Add11~25_combout ),
	.cin(gnd),
	.combout(\Add11~27_combout ),
	.cout());
defparam \Add11~27 .lut_mask = 16'h7FFF;
defparam \Add11~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector119~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[6]~q ),
	.datab(\trk_block:sig_trk_state.s_trk_idle~q ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.cin(gnd),
	.combout(\Selector119~0_combout ),
	.cout());
defparam \Selector119~0 .lut_mask = 16'hEEFF;
defparam \Selector119~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector119~1 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[6]~q ),
	.datab(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datac(\Add10~12_combout ),
	.datad(\shift_in_mmc_seq_value~0_combout ),
	.cin(gnd),
	.combout(\Selector119~1_combout ),
	.cout());
defparam \Selector119~1 .lut_mask = 16'hFAFC;
defparam \Selector119~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector119~2 (
	.dataa(\Selector119~0_combout ),
	.datab(\Selector119~1_combout ),
	.datac(\Equal10~0_combout ),
	.datad(\Equal10~1_combout ),
	.cin(gnd),
	.combout(\Selector119~2_combout ),
	.cout());
defparam \Selector119~2 .lut_mask = 16'hEFFF;
defparam \Selector119~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector122~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector122~0_combout ),
	.cout());
defparam \Selector122~0 .lut_mask = 16'hAAFF;
defparam \Selector122~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~18 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(\sig_req_rsc_shift~54_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add17~18_combout ),
	.cout());
defparam \Add17~18 .lut_mask = 16'hFEFE;
defparam \Add17~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~19 (
	.dataa(\trk_block:sig_mimic_cdv_found~q ),
	.datab(\Add17~1_combout ),
	.datac(\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datad(\sig_dgrb_state.s_track~q ),
	.cin(gnd),
	.combout(\Add17~19_combout ),
	.cout());
defparam \Add17~19 .lut_mask = 16'hFEFF;
defparam \Add17~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~20 (
	.dataa(\Add17~16_combout ),
	.datab(\Add17~18_combout ),
	.datac(\Add17~19_combout ),
	.datad(\trk_block:sig_rsc_drift[7]~q ),
	.cin(gnd),
	.combout(\Add17~20_combout ),
	.cout());
defparam \Add17~20 .lut_mask = 16'hFF7F;
defparam \Add17~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector95~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[6]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector95~0_combout ),
	.cout());
defparam \Selector95~0 .lut_mask = 16'hFEFE;
defparam \Selector95~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~21 (
	.dataa(\Add17~14_combout ),
	.datab(\trk_block:sig_rsc_drift[6]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~21_combout ),
	.cout());
defparam \Add17~21 .lut_mask = 16'hFAFC;
defparam \Add17~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~40 (
	.dataa(\trk_block:sig_rsc_drift[6]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~40_combout ),
	.cout());
defparam \sig_rsc_drift~40 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~40 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector96~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[5]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector96~0_combout ),
	.cout());
defparam \Selector96~0 .lut_mask = 16'hFEFE;
defparam \Selector96~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~22 (
	.dataa(\Add17~12_combout ),
	.datab(\trk_block:sig_rsc_drift[5]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~22_combout ),
	.cout());
defparam \Add17~22 .lut_mask = 16'hFAFC;
defparam \Add17~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~41 (
	.dataa(\trk_block:sig_rsc_drift[5]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~41_combout ),
	.cout());
defparam \sig_rsc_drift~41 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~41 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector69~2 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector69~2_combout ),
	.cout());
defparam \Selector69~2 .lut_mask = 16'hEEEE;
defparam \Selector69~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector97~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[4]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector97~0_combout ),
	.cout());
defparam \Selector97~0 .lut_mask = 16'hFEFE;
defparam \Selector97~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~23 (
	.dataa(\Add17~10_combout ),
	.datab(\trk_block:sig_rsc_drift[4]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~23_combout ),
	.cout());
defparam \Add17~23 .lut_mask = 16'hFAFC;
defparam \Add17~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~42 (
	.dataa(\trk_block:sig_rsc_drift[4]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~42_combout ),
	.cout());
defparam \sig_rsc_drift~42 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~42 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector70~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector70~0_combout ),
	.cout());
defparam \Selector70~0 .lut_mask = 16'hEEEE;
defparam \Selector70~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector98~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[3]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector98~0_combout ),
	.cout());
defparam \Selector98~0 .lut_mask = 16'hFEFE;
defparam \Selector98~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~24 (
	.dataa(\Add17~8_combout ),
	.datab(\trk_block:sig_rsc_drift[3]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~24_combout ),
	.cout());
defparam \Add17~24 .lut_mask = 16'hFAFC;
defparam \Add17~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~43 (
	.dataa(\trk_block:sig_rsc_drift[3]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~43_combout ),
	.cout());
defparam \sig_rsc_drift~43 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~43 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector71~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector71~0_combout ),
	.cout());
defparam \Selector71~0 .lut_mask = 16'hEEEE;
defparam \Selector71~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector99~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[2]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector99~0_combout ),
	.cout());
defparam \Selector99~0 .lut_mask = 16'hFEFE;
defparam \Selector99~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~25 (
	.dataa(\Add17~6_combout ),
	.datab(\trk_block:sig_rsc_drift[2]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~25_combout ),
	.cout());
defparam \Add17~25 .lut_mask = 16'hFAFC;
defparam \Add17~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~44 (
	.dataa(\trk_block:sig_rsc_drift[2]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~44_combout ),
	.cout());
defparam \sig_rsc_drift~44 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~44 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector72~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector72~0_combout ),
	.cout());
defparam \Selector72~0 .lut_mask = 16'hEEEE;
defparam \Selector72~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector100~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_rsc_drift[1]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector100~0_combout ),
	.cout());
defparam \Selector100~0 .lut_mask = 16'hFEFE;
defparam \Selector100~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~26 (
	.dataa(\Add17~4_combout ),
	.datab(\trk_block:sig_rsc_drift[1]~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\sig_req_rsc_shift~54_combout ),
	.cin(gnd),
	.combout(\Add17~26_combout ),
	.cout());
defparam \Add17~26 .lut_mask = 16'hFAFC;
defparam \Add17~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_drift~45 (
	.dataa(\trk_block:sig_rsc_drift[1]~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_rsc_drift~45_combout ),
	.cout());
defparam \sig_rsc_drift~45 .lut_mask = 16'hEEEE;
defparam \sig_rsc_drift~45 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector73~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector73~0_combout ),
	.cout());
defparam \Selector73~0 .lut_mask = 16'hEEEE;
defparam \Selector73~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~27 (
	.dataa(\Add17~18_combout ),
	.datab(\Add17~19_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_rsc_drift[0]~q ),
	.cin(gnd),
	.combout(\Add17~27_combout ),
	.cout());
defparam \Add17~27 .lut_mask = 16'h5533;
defparam \Add17~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_test_dq_expired~6 (
	.dataa(\rsc_block:sig_count[0]~q ),
	.datab(\Equal7~1_combout ),
	.datac(\sig_dimm_driving_dq~q ),
	.datad(\rsc_proc~1_combout ),
	.cin(gnd),
	.combout(\sig_test_dq_expired~6_combout ),
	.cout());
defparam \sig_test_dq_expired~6 .lut_mask = 16'hEFFF;
defparam \sig_test_dq_expired~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal8~0 (
	.dataa(\tp_match_block:sig_rdata_current_pin[13]~q ),
	.datab(\tp_match_block:sig_rdata_current_pin[12]~q ),
	.datac(\tp_match_block:sig_rdata_current_pin[11]~q ),
	.datad(\tp_match_block:sig_rdata_current_pin[10]~q ),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
defparam \Equal8~0 .lut_mask = 16'hEFFF;
defparam \Equal8~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~434 (
	.dataa(\sig_cdvw_state.current_window_centre[5]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~434_combout ),
	.cout());
defparam \v_cdvw_state~434 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~434 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~435 (
	.dataa(\sig_cdvw_state.current_window_centre[4]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~435_combout ),
	.cout());
defparam \v_cdvw_state~435 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~435 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~436 (
	.dataa(\sig_cdvw_state.current_window_centre[3]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~436_combout ),
	.cout());
defparam \v_cdvw_state~436 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~436 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~437 (
	.dataa(\sig_cdvw_state.current_window_centre[2]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~437_combout ),
	.cout());
defparam \v_cdvw_state~437 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~437 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~438 (
	.dataa(\sig_cdvw_state.current_window_centre[1]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~438_combout ),
	.cout());
defparam \v_cdvw_state~438 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~438 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~441 (
	.dataa(\sig_cdvw_state.current_bit[2]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~441_combout ),
	.cout());
defparam \v_cdvw_state~441 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~441 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~442 (
	.dataa(\sig_cdvw_state.current_bit[5]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~442_combout ),
	.cout());
defparam \v_cdvw_state~442 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~442 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~447 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.invalid_phase_seen~q ),
	.datac(\sig_cdvw_state.status.calculating~q ),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~447_combout ),
	.cout());
defparam \v_cdvw_state~447 .lut_mask = 16'hFFFE;
defparam \v_cdvw_state~447 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~450 (
	.dataa(\sig_cdvw_state.largest_window_size[5]~q ),
	.datab(\sig_cdvw_state.largest_window_size[2]~q ),
	.datac(\sig_cdvw_state.current_window_size[2]~q ),
	.datad(\sig_cdvw_state.current_window_size[5]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~450_combout ),
	.cout());
defparam \v_cdvw_state~450 .lut_mask = 16'h6996;
defparam \v_cdvw_state~450 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\Selector50~0_combout ),
	.cout());
defparam \Selector50~0 .lut_mask = 16'hEEFF;
defparam \Selector50~0 .sum_lutc_input = "datac";

dffeas \tp_match_block:sig_rdata_valid_2t (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_valid_1t~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_valid_2t~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_valid_2t .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_valid_2t .power_up = "low";

cycloneiii_lcell_comb \trk_block:sig_mimic_cdv[0]~1 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_cdvw_state.status.valid_result~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\trk_block:sig_mimic_cdv[0]~1_combout ),
	.cout());
defparam \trk_block:sig_mimic_cdv[0]~1 .lut_mask = 16'hFEFE;
defparam \trk_block:sig_mimic_cdv[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector35~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\single_bit_cal~q ),
	.cin(gnd),
	.combout(\Selector35~0_combout ),
	.cout());
defparam \Selector35~0 .lut_mask = 16'hAAFF;
defparam \Selector35~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~0 (
	.dataa(\sig_dq_pin_ctr[2]~q ),
	.datab(q_b_25),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_9),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~1 (
	.dataa(q_b_13),
	.datab(\sig_dq_pin_ctr[2]~q ),
	.datac(\Mux1~0_combout ),
	.datad(q_b_29),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~0 (
	.dataa(\sig_dq_pin_ctr[1]~q ),
	.datab(q_b_17),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_1),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~1 (
	.dataa(q_b_3),
	.datab(\sig_dq_pin_ctr[1]~q ),
	.datac(\Mux0~0_combout ),
	.datad(q_b_19),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~18 (
	.dataa(\sig_cdvw_state.current_window_centre[0]~q ),
	.datab(\sig_cdvw_state.current_window_centre[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[5]~18_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~18 .lut_mask = 16'hEEEE;
defparam \sig_cdvw_state.current_window_centre[5]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~19 (
	.dataa(\sig_cdvw_state.current_window_centre[4]~q ),
	.datab(\sig_cdvw_state.current_window_centre[3]~q ),
	.datac(\sig_cdvw_state.current_window_centre[2]~q ),
	.datad(\sig_cdvw_state.current_window_centre[1]~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[5]~19_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~19 .lut_mask = 16'hFFFE;
defparam \sig_cdvw_state.current_window_centre[5]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~20 (
	.dataa(\sig_cdvw_state.current_window_centre[5]~18_combout ),
	.datab(\sig_cdvw_state.current_window_centre[5]~19_combout ),
	.datac(\find_centre_of_largest_data_valid_window~6_combout ),
	.datad(\v_cdvw_state~430_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[5]~20_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~20 .lut_mask = 16'hEFFF;
defparam \sig_cdvw_state.current_window_centre[5]~20 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.window_centre_update (
	.clk(clk),
	.d(\v_cdvw_state~465_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.window_centre_update~q ),
	.prn(vcc));
defparam \sig_cdvw_state.window_centre_update .is_wysiwyg = "true";
defparam \sig_cdvw_state.window_centre_update .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~21 (
	.dataa(\sig_cdvw_state.window_centre_update~q ),
	.datab(gnd),
	.datac(\sig_cdvw_state.found_a_good_edge~q ),
	.datad(\sig_cdvw_state.last_bit_value~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[5]~21_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~21 .lut_mask = 16'hAFFF;
defparam \sig_cdvw_state.current_window_centre[5]~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_centre[5]~22 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.working_window[0]~q ),
	.datac(\sig_cdvw_state.current_window_centre[5]~21_combout ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_centre[5]~22_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_centre[5]~22 .lut_mask = 16'hFF7F;
defparam \sig_cdvw_state.current_window_centre[5]~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[0]~19 (
	.dataa(\sig_cdvw_state.working_window[0]~q ),
	.datab(\sig_cdvw_state.last_bit_value~q ),
	.datac(\sig_cdvw_state.found_a_good_edge~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~19_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_size[0]~19 .lut_mask = 16'h6FFF;
defparam \sig_cdvw_state.current_window_size[0]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~464 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\sig_cdvw_state.found_a_good_edge~q ),
	.datac(\sig_cdvw_state.last_bit_value~q ),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~464_combout ),
	.cout());
defparam \v_cdvw_state~464 .lut_mask = 16'hFEFF;
defparam \v_cdvw_state~464 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~465 (
	.dataa(\v_cdvw_state~464_combout ),
	.datab(\find_centre_of_largest_data_valid_window~7_combout ),
	.datac(\sig_cdvw_state.window_centre_update~q ),
	.datad(\v_cdvw_state~430_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~465_combout ),
	.cout());
defparam \v_cdvw_state~465 .lut_mask = 16'hFF7B;
defparam \v_cdvw_state~465 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_last_state.s_trk_mimic_sample (
	.clk(clk),
	.d(\sig_trk_last_state~31_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_mimic_sample~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_mimic_sample .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_mimic_sample .power_up = "low";

cycloneiii_lcell_comb \sig_trk_last_state~31 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_last_state~31_combout ),
	.cout());
defparam \sig_trk_last_state~31 .lut_mask = 16'hEEEE;
defparam \sig_trk_last_state~31 .sum_lutc_input = "datac";

dffeas sig_trk_cdvw_phase(
	.clk(clk),
	.d(\sig_trk_cdvw_phase~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_phase~q ),
	.prn(vcc));
defparam sig_trk_cdvw_phase.is_wysiwyg = "true";
defparam sig_trk_cdvw_phase.power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~528 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_cdvw_phase~q ),
	.datac(\sig_rsc_cdvw_phase~q ),
	.datad(\WideOr11~2_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~528_combout ),
	.cout());
defparam \v_cdvw_state~528 .lut_mask = 16'hFEFF;
defparam \v_cdvw_state~528 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~529 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\v_cdvw_state~528_combout ),
	.datac(gnd),
	.datad(\sig_cdvw_state.working_window[12]~4_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~529_combout ),
	.cout());
defparam \v_cdvw_state~529 .lut_mask = 16'hEEFF;
defparam \v_cdvw_state~529 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_cdvw_phase~1 (
	.dataa(\trk_block:sig_mmc_seq_done_1t~q ),
	.datab(mimic_value_captured),
	.datac(gnd),
	.datad(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.cin(gnd),
	.combout(\sig_trk_cdvw_phase~1_combout ),
	.cout());
defparam \sig_trk_cdvw_phase~1 .lut_mask = 16'hEEFF;
defparam \sig_trk_cdvw_phase~1 .sum_lutc_input = "datac";

dffeas \rsc_block:rsc_proc:v_phase_works (
	.clk(clk),
	.d(\Selector66~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:rsc_proc:v_phase_works~q ),
	.prn(vcc));
defparam \rsc_block:rsc_proc:v_phase_works .is_wysiwyg = "true";
defparam \rsc_block:rsc_proc:v_phase_works .power_up = "low";

cycloneiii_lcell_comb \rsc_proc~3 (
	.dataa(\rsc_block:sig_curr_byte_ln_dis~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_mtp_match~q ),
	.cin(gnd),
	.combout(\rsc_proc~3_combout ),
	.cout());
defparam \rsc_proc~3 .lut_mask = 16'hAAFF;
defparam \rsc_proc~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_cdvw_phase~5 (
	.dataa(\rsc_block:sig_chkd_all_dq_pins~q ),
	.datab(\rsc_block:rsc_proc:v_phase_works~q ),
	.datac(\sig_dimm_driving_dq~q ),
	.datad(\rsc_proc~3_combout ),
	.cin(gnd),
	.combout(\sig_rsc_cdvw_phase~5_combout ),
	.cout());
defparam \sig_rsc_cdvw_phase~5 .lut_mask = 16'hEFFF;
defparam \sig_rsc_cdvw_phase~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector66~0 (
	.dataa(\sig_dimm_driving_dq~q ),
	.datab(\rsc_block:sig_test_dq_expired~q ),
	.datac(\rsc_proc~3_combout ),
	.datad(\rsc_block:sig_count[6]~5_combout ),
	.cin(gnd),
	.combout(\Selector66~0_combout ),
	.cout());
defparam \Selector66~0 .lut_mask = 16'hBFFF;
defparam \Selector66~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector66~1 (
	.dataa(\rsc_block:rsc_proc:v_phase_works~q ),
	.datab(\Selector66~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\Selector66~1_combout ),
	.cout());
defparam \Selector66~1 .lut_mask = 16'hFEFF;
defparam \Selector66~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~68 (
	.dataa(\LessThan10~1_combout ),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(\Add16~12_combout ),
	.datad(\Add18~12_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~68_combout ),
	.cout());
defparam \sig_req_rsc_shift~68 .lut_mask = 16'hF7D5;
defparam \sig_req_rsc_shift~68 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector42~3 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(\Selector42~2_combout ),
	.datad(\sig_cdvw_state.largest_window_centre[4]~q ),
	.cin(gnd),
	.combout(\Selector42~3_combout ),
	.cout());
defparam \Selector42~3 .lut_mask = 16'hFFFD;
defparam \Selector42~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~28 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~12_combout ),
	.cin(gnd),
	.combout(\Add11~28_combout ),
	.cout());
defparam \Add11~28 .lut_mask = 16'hFFFE;
defparam \Add11~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~29 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~23_combout ),
	.cin(gnd),
	.combout(\Add11~29_combout ),
	.cout());
defparam \Add11~29 .lut_mask = 16'hFFFE;
defparam \Add11~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~30 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~21_combout ),
	.cin(gnd),
	.combout(\Add11~30_combout ),
	.cout());
defparam \Add11~30 .lut_mask = 16'hFFFE;
defparam \Add11~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~31 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~19_combout ),
	.cin(gnd),
	.combout(\Add11~31_combout ),
	.cout());
defparam \Add11~31 .lut_mask = 16'hFFFE;
defparam \Add11~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~32 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~17_combout ),
	.cin(gnd),
	.combout(\Add11~32_combout ),
	.cout());
defparam \Add11~32 .lut_mask = 16'hFFFE;
defparam \Add11~32 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add11~33 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_mimic_cdv_found~q ),
	.datad(\Add11~15_combout ),
	.cin(gnd),
	.combout(\Add11~33_combout ),
	.cout());
defparam \Add11~33 .lut_mask = 16'hFFFE;
defparam \Add11~33 .sum_lutc_input = "datac";

dffeas \sig_doing_rd[0] (
	.clk(clk),
	.d(\Selector175~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_doing_rd_0),
	.prn(vcc));
defparam \sig_doing_rd[0] .is_wysiwyg = "true";
defparam \sig_doing_rd[0] .power_up = "low";

dffeas \sig_doing_rd[1] (
	.clk(clk),
	.d(\Selector175~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_doing_rd_1),
	.prn(vcc));
defparam \sig_doing_rd[1] .is_wysiwyg = "true";
defparam \sig_doing_rd[1] .power_up = "low";

dffeas dgrb_ac_access_req(
	.clk(clk),
	.d(\dimm_driving_dq_proc~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ac_access_req1),
	.prn(vcc));
defparam dgrb_ac_access_req.is_wysiwyg = "true";
defparam dgrb_ac_access_req.power_up = "low";

dffeas \sig_addr_cmd[0].cs_n[0] (
	.clk(clk),
	.d(\Selector165~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0cs_n0),
	.prn(vcc));
defparam \sig_addr_cmd[0].cs_n[0] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cs_n[0] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[2] (
	.clk(clk),
	.d(\Selector141~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr2),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[2] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[2] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[3] (
	.clk(clk),
	.d(\Selector140~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr3),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[3] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[3] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[4] (
	.clk(clk),
	.d(\Selector139~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr4),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[4] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[4] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[5] (
	.clk(clk),
	.d(\Selector138~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr5),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[5] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[5] .power_up = "low";

dffeas \sig_addr_cmd[0].cas_n (
	.clk(clk),
	.d(\sig_addr_cmd[0].cas_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0cas_n),
	.prn(vcc));
defparam \sig_addr_cmd[0].cas_n .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cas_n .power_up = "low";

dffeas \wd_lat[0] (
	.clk(clk),
	.d(\wd_lat[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_0),
	.prn(vcc));
defparam \wd_lat[0] .is_wysiwyg = "true";
defparam \wd_lat[0] .power_up = "low";

dffeas \wd_lat[1] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_1),
	.prn(vcc));
defparam \wd_lat[1] .is_wysiwyg = "true";
defparam \wd_lat[1] .power_up = "low";

dffeas \wd_lat[4] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_4),
	.prn(vcc));
defparam \wd_lat[4] .is_wysiwyg = "true";
defparam \wd_lat[4] .power_up = "low";

dffeas \wd_lat[3] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_3),
	.prn(vcc));
defparam \wd_lat[3] .is_wysiwyg = "true";
defparam \wd_lat[3] .power_up = "low";

dffeas \wd_lat[2] (
	.clk(clk),
	.d(\wd_lat[2]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_2),
	.prn(vcc));
defparam \wd_lat[2] .is_wysiwyg = "true";
defparam \wd_lat[2] .power_up = "low";

dffeas seq_rdata_valid_lat_dec(
	.clk(clk),
	.d(\seq_rdata_valid_lat_dec~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_lat_dec1),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec.power_up = "low";

dffeas seq_pll_inc_dec_n(
	.clk(clk),
	.d(\seq_pll_inc_dec_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_inc_dec_n1),
	.prn(vcc));
defparam seq_pll_inc_dec_n.is_wysiwyg = "true";
defparam seq_pll_inc_dec_n.power_up = "low";

dffeas seq_pll_start_reconfig(
	.clk(clk),
	.d(\seq_pll_start_reconfig~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_start_reconfig1),
	.prn(vcc));
defparam seq_pll_start_reconfig.is_wysiwyg = "true";
defparam seq_pll_start_reconfig.power_up = "low";

dffeas \dgrb_ctrl.command_done (
	.clk(clk),
	.d(\ac_handshake_proc~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_done),
	.prn(vcc));
defparam \dgrb_ctrl.command_done .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_done .power_up = "low";

dffeas \seq_pll_select[2] (
	.clk(clk),
	.d(\seq_pll_select~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_2),
	.prn(vcc));
defparam \seq_pll_select[2] .is_wysiwyg = "true";
defparam \seq_pll_select[2] .power_up = "low";

dffeas \seq_pll_select[0] (
	.clk(clk),
	.d(\seq_pll_select~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_0),
	.prn(vcc));
defparam \seq_pll_select[0] .is_wysiwyg = "true";
defparam \seq_pll_select[0] .power_up = "low";

dffeas \dgrb_ctrl.command_result[5] (
	.clk(clk),
	.d(\dgrb_ctrl~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_5),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[5] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[5] .power_up = "low";

dffeas \dgrb_ctrl.command_result[4] (
	.clk(clk),
	.d(\dgrb_ctrl~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_4),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[4] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[4] .power_up = "low";

dffeas \dgrb_ctrl.command_result[3] (
	.clk(clk),
	.d(\dgrb_ctrl~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_3),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[3] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[3] .power_up = "low";

dffeas \dgrb_ctrl.command_result[2] (
	.clk(clk),
	.d(\dgrb_ctrl~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_2),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[2] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[2] .power_up = "low";

dffeas \dgrb_ctrl.command_result[1] (
	.clk(clk),
	.d(\dgrb_ctrl~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_1),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[1] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[1] .power_up = "low";

dffeas \dgrb_ctrl.command_result[0] (
	.clk(clk),
	.d(\dgrb_ctrl~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_0),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[0] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[0] .power_up = "low";

dffeas seq_mmc_start(
	.clk(clk),
	.d(\seq_mmc_start~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_mmc_start1),
	.prn(vcc));
defparam seq_mmc_start.is_wysiwyg = "true";
defparam seq_mmc_start.power_up = "low";

cycloneiii_lcell_comb \Add23~6 (
	.dataa(\ac_block:sig_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~5 ),
	.combout(\Add23~6_combout ),
	.cout(\Add23~7 ));
defparam \Add23~6 .lut_mask = 16'h5A5F;
defparam \Add23~6 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add23~8 (
	.dataa(\ac_block:sig_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~7 ),
	.combout(\Add23~8_combout ),
	.cout(\Add23~9 ));
defparam \Add23~8 .lut_mask = 16'h5AAF;
defparam \Add23~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add23~10 (
	.dataa(\ac_block:sig_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add23~9 ),
	.combout(\Add23~10_combout ),
	.cout(\Add23~11 ));
defparam \Add23~10 .lut_mask = 16'h5A5F;
defparam \Add23~10 .sum_lutc_input = "cin";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~237 (
	.dataa(q_b_0),
	.datab(q_b_8),
	.datac(gnd),
	.datad(rdata_valid[0]),
	.cin(gnd),
	.combout(\sig_dgrb_state~237_combout ),
	.cout());
defparam \sig_dgrb_state~237 .lut_mask = 16'hEEFF;
defparam \sig_dgrb_state~237 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~261 (
	.dataa(\sig_dimm_driving_dq~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\sig_dgrb_state~261_combout ),
	.cout());
defparam \sig_dgrb_state~261 .lut_mask = 16'hAAFF;
defparam \sig_dgrb_state~261 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~262 (
	.dataa(WideOr1),
	.datab(\sig_dgrb_state.s_release_admin~q ),
	.datac(\sig_dgrb_state~261_combout ),
	.datad(\sig_dgrb_state.s_wait_admin~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~262_combout ),
	.cout());
defparam \sig_dgrb_state~262 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~262 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~264 (
	.dataa(last_states_adv_wr_lat),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~264_combout ),
	.cout());
defparam \sig_dgrb_state~264 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~264 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~281 (
	.dataa(curr_cmdcmd_idle),
	.datab(\sig_dgrb_state.s_release_admin~q ),
	.datac(\sig_dgrb_state.s_idle~q ),
	.datad(\sig_dgrb_state~257_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~281_combout ),
	.cout());
defparam \sig_dgrb_state~281 .lut_mask = 16'hF7FF;
defparam \sig_dgrb_state~281 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_adv_wd_lat (
	.clk(clk),
	.d(\sig_dgrb_state~264_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_adv_wd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_wd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_wd_lat .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~268 (
	.dataa(ac_muxctrl_broadcast_rcommand_req),
	.datab(gnd),
	.datac(WideOr1),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~268_combout ),
	.cout());
defparam \sig_dgrb_state~268 .lut_mask = 16'hAFFF;
defparam \sig_dgrb_state~268 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~269 (
	.dataa(\sig_dgrb_state.s_adv_rd_lat~q ),
	.datab(\sig_dgrb_state~267_combout ),
	.datac(gnd),
	.datad(\sig_dgrb_state~268_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~269_combout ),
	.cout());
defparam \sig_dgrb_state~269 .lut_mask = 16'hEEFF;
defparam \sig_dgrb_state~269 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~259 (
	.dataa(last_states_rrp_reset),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~259_combout ),
	.cout());
defparam \sig_dgrb_state~259 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~259 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_reset_cdvw (
	.clk(clk),
	.d(\sig_dgrb_state~259_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_reset_cdvw~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_reset_cdvw .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_reset_cdvw .power_up = "low";

cycloneiii_lcell_comb \sig_rsc_req~28 (
	.dataa(\sig_rsc_ack~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_reset_cdvw~q ),
	.cin(gnd),
	.combout(\sig_rsc_req~28_combout ),
	.cout());
defparam \sig_rsc_req~28 .lut_mask = 16'hFF55;
defparam \sig_rsc_req~28 .sum_lutc_input = "datac";

dffeas \sig_rsc_req.s_rsc_reset_cdvw (
	.clk(clk),
	.d(\sig_rsc_req~28_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_reset_cdvw .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_reset_cdvw .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_idle (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_idle .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_idle .power_up = "low";

cycloneiii_lcell_comb \Selector54~0 (
	.dataa(\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.datab(gnd),
	.datac(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datad(\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.cin(gnd),
	.combout(\Selector54~0_combout ),
	.cout());
defparam \Selector54~0 .lut_mask = 16'hAFFF;
defparam \Selector54~0 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_reset_cdvw (
	.clk(clk),
	.d(\Selector54~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_reset_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_reset_cdvw .power_up = "low";

cycloneiii_lcell_comb \Selector37~0 (
	.dataa(\Selector35~0_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(\sig_dq_pin_ctr[1]~q ),
	.datad(\sig_dq_pin_ctr[0]~q ),
	.cin(gnd),
	.combout(\Selector37~0_combout ),
	.cout());
defparam \Selector37~0 .lut_mask = 16'hEFFE;
defparam \Selector37~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr12~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.cin(gnd),
	.combout(\WideOr12~0_combout ),
	.cout());
defparam \WideOr12~0 .lut_mask = 16'hAAFF;
defparam \WideOr12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dq_pin_ctr[3]~16 (
	.dataa(\rsc_block:sig_chkd_all_dq_pins~q ),
	.datab(\WideOr12~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Selector51~0_combout ),
	.cin(gnd),
	.combout(\sig_dq_pin_ctr[3]~16_combout ),
	.cout());
defparam \sig_dq_pin_ctr[3]~16 .lut_mask = 16'hF737;
defparam \sig_dq_pin_ctr[3]~16 .sum_lutc_input = "datac";

dffeas \sig_dq_pin_ctr[1] (
	.clk(clk),
	.d(\Selector37~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dq_pin_ctr[3]~16_combout ),
	.q(\sig_dq_pin_ctr[1]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[1] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[1] .power_up = "low";

cycloneiii_lcell_comb \Equal4~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sig_dq_pin_ctr[1]~q ),
	.datad(\sig_dq_pin_ctr[0]~q ),
	.cin(gnd),
	.combout(\Equal4~2_combout ),
	.cout());
defparam \Equal4~2 .lut_mask = 16'h0FFF;
defparam \Equal4~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector36~0 (
	.dataa(\Selector35~0_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(\sig_dq_pin_ctr[2]~q ),
	.datad(\Equal4~2_combout ),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hEFFE;
defparam \Selector36~0 .sum_lutc_input = "datac";

dffeas \sig_dq_pin_ctr[2] (
	.clk(clk),
	.d(\Selector36~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dq_pin_ctr[3]~16_combout ),
	.q(\sig_dq_pin_ctr[2]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[2] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[2] .power_up = "low";

cycloneiii_lcell_comb \Equal4~1 (
	.dataa(gnd),
	.datab(\sig_dq_pin_ctr[2]~q ),
	.datac(\sig_dq_pin_ctr[1]~q ),
	.datad(\sig_dq_pin_ctr[0]~q ),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
defparam \Equal4~1 .lut_mask = 16'h3FFF;
defparam \Equal4~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector35~1 (
	.dataa(\Selector35~0_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(\Equal4~1_combout ),
	.cin(gnd),
	.combout(\Selector35~1_combout ),
	.cout());
defparam \Selector35~1 .lut_mask = 16'hEFFE;
defparam \Selector35~1 .sum_lutc_input = "datac";

dffeas \sig_dq_pin_ctr[3] (
	.clk(clk),
	.d(\Selector35~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dq_pin_ctr[3]~16_combout ),
	.q(\sig_dq_pin_ctr[3]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[3] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[3] .power_up = "low";

cycloneiii_lcell_comb \Mux0~2 (
	.dataa(\sig_dq_pin_ctr[1]~q ),
	.datab(q_b_20),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_4),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFDE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~3 (
	.dataa(q_b_6),
	.datab(\sig_dq_pin_ctr[1]~q ),
	.datac(\Mux0~2_combout ),
	.datad(q_b_22),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFBE;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~4 (
	.dataa(\sig_dq_pin_ctr[1]~q ),
	.datab(q_b_16),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_0),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hFFDE;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~5 (
	.dataa(q_b_2),
	.datab(\sig_dq_pin_ctr[1]~q ),
	.datac(\Mux0~4_combout ),
	.datad(q_b_18),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hFFBE;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~6 (
	.dataa(\sig_dq_pin_ctr[0]~q ),
	.datab(\Mux0~3_combout ),
	.datac(\sig_dq_pin_ctr[2]~q ),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
defparam \Mux0~6 .lut_mask = 16'hFFDE;
defparam \Mux0~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~7 (
	.dataa(\sig_dq_pin_ctr[1]~q ),
	.datab(q_b_21),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_5),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
defparam \Mux0~7 .lut_mask = 16'hFFDE;
defparam \Mux0~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~8 (
	.dataa(q_b_7),
	.datab(\sig_dq_pin_ctr[1]~q ),
	.datac(\Mux0~7_combout ),
	.datad(q_b_23),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
defparam \Mux0~8 .lut_mask = 16'hFFBE;
defparam \Mux0~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux0~9 (
	.dataa(\Mux0~1_combout ),
	.datab(\sig_dq_pin_ctr[0]~q ),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~8_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
defparam \Mux0~9 .lut_mask = 16'hFFBE;
defparam \Mux0~9 .sum_lutc_input = "datac";

dffeas \tp_match_block:sig_rdata_current_pin[14] (
	.clk(clk),
	.d(\Mux0~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[14] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[14] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[13] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[13]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[13] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[13] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[11] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[13]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[11]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[11] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[11] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[9] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[11]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[9]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[9] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[9] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[12] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[12]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[12] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[12] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[10] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[12]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[10]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[10] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[10] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[8] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[10]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[8]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[8] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[8] .power_up = "low";

cycloneiii_lcell_comb \Equal8~1 (
	.dataa(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.datab(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.datac(\tp_match_block:sig_rdata_current_pin[9]~q ),
	.datad(\tp_match_block:sig_rdata_current_pin[8]~q ),
	.cin(gnd),
	.combout(\Equal8~1_combout ),
	.cout());
defparam \Equal8~1 .lut_mask = 16'h7FFF;
defparam \Equal8~1 .sum_lutc_input = "datac";

dffeas \tp_match_block:sig_rdata_current_pin[6] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[8]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[6]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[6] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[6] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[7] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[9]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[7]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[7] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[7] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[5] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[7]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[5]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[5] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[5] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[4] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[6]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[4]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[4] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[4] .power_up = "low";

cycloneiii_lcell_comb \Equal8~2 (
	.dataa(\tp_match_block:sig_rdata_current_pin[7]~q ),
	.datab(\tp_match_block:sig_rdata_current_pin[6]~q ),
	.datac(\tp_match_block:sig_rdata_current_pin[5]~q ),
	.datad(\tp_match_block:sig_rdata_current_pin[4]~q ),
	.cin(gnd),
	.combout(\Equal8~2_combout ),
	.cout());
defparam \Equal8~2 .lut_mask = 16'hFFFE;
defparam \Equal8~2 .sum_lutc_input = "datac";

dffeas \tp_match_block:sig_rdata_current_pin[2] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[2]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[2] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[2] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[0] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[0]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[0] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[0] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[3] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[3]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[3] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[3] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[1] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[1]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[1] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[1] .power_up = "low";

cycloneiii_lcell_comb \Equal8~3 (
	.dataa(\tp_match_block:sig_rdata_current_pin[2]~q ),
	.datab(\tp_match_block:sig_rdata_current_pin[0]~q ),
	.datac(\tp_match_block:sig_rdata_current_pin[3]~q ),
	.datad(\tp_match_block:sig_rdata_current_pin[1]~q ),
	.cin(gnd),
	.combout(\Equal8~3_combout ),
	.cout());
defparam \Equal8~3 .lut_mask = 16'hEFFF;
defparam \Equal8~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal8~4 (
	.dataa(\Equal8~0_combout ),
	.datab(\Equal8~1_combout ),
	.datac(\Equal8~2_combout ),
	.datad(\Equal8~3_combout ),
	.cin(gnd),
	.combout(\Equal8~4_combout ),
	.cout());
defparam \Equal8~4 .lut_mask = 16'hFFFE;
defparam \Equal8~4 .sum_lutc_input = "datac";

dffeas sig_mtp_match(
	.clk(clk),
	.d(\Equal8~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_mtp_match~q ),
	.prn(vcc));
defparam sig_mtp_match.is_wysiwyg = "true";
defparam sig_mtp_match.power_up = "low";

dffeas \rsc_block:sig_curr_byte_ln_dis (
	.clk(clk),
	.d(seq_ac_add_1t_ac_lat_internal),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_curr_byte_ln_dis~q ),
	.prn(vcc));
defparam \rsc_block:sig_curr_byte_ln_dis .is_wysiwyg = "true";
defparam \rsc_block:sig_curr_byte_ln_dis .power_up = "low";

cycloneiii_lcell_comb \rsc_proc~1 (
	.dataa(\rsc_block:sig_test_dq_expired~q ),
	.datab(\sig_mtp_match~q ),
	.datac(gnd),
	.datad(\rsc_block:sig_curr_byte_ln_dis~q ),
	.cin(gnd),
	.combout(\rsc_proc~1_combout ),
	.cout());
defparam \rsc_proc~1 .lut_mask = 16'hEEFF;
defparam \rsc_proc~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector51~0 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datab(\rsc_proc~1_combout ),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\Selector51~0_combout ),
	.cout());
defparam \Selector51~0 .lut_mask = 16'hEEFF;
defparam \Selector51~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector52~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(\Selector52~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Selector51~0_combout ),
	.cin(gnd),
	.combout(\Selector52~1_combout ),
	.cout());
defparam \Selector52~1 .lut_mask = 16'hFEFF;
defparam \Selector52~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_test_dq (
	.clk(clk),
	.d(\Selector52~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_test_dq .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_test_dq .power_up = "low";

cycloneiii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~0 (
	.dataa(\Add9~16_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.cout());
defparam \rsc_block:sig_num_phase_shifts[2]~0 .lut_mask = 16'hAAFF;
defparam \rsc_block:sig_num_phase_shifts[2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~0 (
	.dataa(\sig_dq_pin_ctr[3]~q ),
	.datab(\sig_dq_pin_ctr[2]~q ),
	.datac(\sig_dq_pin_ctr[1]~q ),
	.datad(\sig_dq_pin_ctr[0]~q ),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h7FFF;
defparam \Equal4~0 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_chkd_all_dq_pins (
	.clk(clk),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_chkd_all_dq_pins~q ),
	.prn(vcc));
defparam \rsc_block:sig_chkd_all_dq_pins .is_wysiwyg = "true";
defparam \rsc_block:sig_chkd_all_dq_pins .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_test_dq (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_test_dq .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_test_dq .power_up = "low";

cycloneiii_lcell_comb \Selector51~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(\rsc_proc~1_combout ),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\Selector51~1_combout ),
	.cout());
defparam \Selector51~1 .lut_mask = 16'hFEFF;
defparam \Selector51~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector48~1 (
	.dataa(\Selector48~0_combout ),
	.datab(\Equal6~1_combout ),
	.datac(\rsc_block:sig_chkd_all_dq_pins~q ),
	.datad(\Selector51~1_combout ),
	.cin(gnd),
	.combout(\Selector48~1_combout ),
	.cout());
defparam \Selector48~1 .lut_mask = 16'hFFFE;
defparam \Selector48~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_next_phase (
	.clk(clk),
	.d(\Selector48~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_next_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_next_phase .power_up = "low";

cycloneiii_lcell_comb \Add5~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.cin(gnd),
	.combout(\Add5~3_combout ),
	.cout());
defparam \Add5~3 .lut_mask = 16'h0FFF;
defparam \Add5~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~9 (
	.dataa(\Add5~1_combout ),
	.datab(\Add5~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add5~9_combout ),
	.cout(\Add5~10 ));
defparam \Add5~9 .lut_mask = 16'h66EE;
defparam \Add5~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~26 (
	.dataa(\Add9~0_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~9_combout ),
	.cin(gnd),
	.combout(\Add5~26_combout ),
	.cout());
defparam \Add5~26 .lut_mask = 16'h47FF;
defparam \Add5~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~1 (
	.dataa(\Equal6~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.cout());
defparam \rsc_block:sig_num_phase_shifts[2]~1 .lut_mask = 16'hFEFE;
defparam \rsc_block:sig_num_phase_shifts[2]~1 .sum_lutc_input = "datac";

dffeas \phs_shft_busy_reg:phs_shft_busy_1r (
	.clk(clk),
	.d(phs_shft_busy),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phs_shft_busy_reg:phs_shft_busy_1r~q ),
	.prn(vcc));
defparam \phs_shft_busy_reg:phs_shft_busy_1r .is_wysiwyg = "true";
defparam \phs_shft_busy_reg:phs_shft_busy_1r .power_up = "low";

dffeas \phs_shft_busy_reg:phs_shft_busy_2r (
	.clk(clk),
	.d(\phs_shft_busy_reg:phs_shft_busy_1r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.prn(vcc));
defparam \phs_shft_busy_reg:phs_shft_busy_2r .is_wysiwyg = "true";
defparam \phs_shft_busy_reg:phs_shft_busy_2r .power_up = "low";

dffeas sig_phs_shft_busy(
	.clk(clk),
	.d(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_busy~q ),
	.prn(vcc));
defparam sig_phs_shft_busy.is_wysiwyg = "true";
defparam sig_phs_shft_busy.power_up = "low";

dffeas sig_phs_shft_busy_1t(
	.clk(clk),
	.d(\sig_phs_shft_busy~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_busy_1t~q ),
	.prn(vcc));
defparam sig_phs_shft_busy_1t.is_wysiwyg = "true";
defparam sig_phs_shft_busy_1t.power_up = "low";

cycloneiii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~2 (
	.dataa(\sig_phs_shft_busy~q ),
	.datab(\sig_phs_shft_busy_1t~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~2_combout ),
	.cout());
defparam \rsc_block:sig_num_phase_shifts[2]~2 .lut_mask = 16'hDFD5;
defparam \rsc_block:sig_num_phase_shifts[2]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~3 (
	.dataa(\sig_phs_shft_end~q ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~2_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datad(\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~3_combout ),
	.cout());
defparam \rsc_block:sig_num_phase_shifts[2]~3 .lut_mask = 16'hEFFE;
defparam \rsc_block:sig_num_phase_shifts[2]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~4 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(\Selector53~0_combout ),
	.datac(\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datad(\rsc_block:sig_num_phase_shifts[2]~3_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.cout());
defparam \rsc_block:sig_num_phase_shifts[2]~4 .lut_mask = 16'hDF8F;
defparam \rsc_block:sig_num_phase_shifts[2]~4 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_num_phase_shifts[0] (
	.clk(clk),
	.d(\Add5~26_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[0]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[0] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[0] .power_up = "low";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r (
	.clk(clk),
	.d(mmc_seq_done),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r .power_up = "low";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r .power_up = "low";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r .power_up = "low";

dffeas \trk_block:sig_mmc_seq_done_1t (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_mmc_seq_done_1t~q ),
	.prn(vcc));
defparam \trk_block:sig_mmc_seq_done_1t .is_wysiwyg = "true";
defparam \trk_block:sig_mmc_seq_done_1t .power_up = "low";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[2]~0 (
	.dataa(\Add10~4_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[2]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[2]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[2]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[2]~0 .sum_lutc_input = "datac";

dffeas \ctrl_dgrb_r.command.cmd_tr_due (
	.clk(clk),
	.d(Selector57),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_tr_due~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_tr_due .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_tr_due .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~241 (
	.dataa(\sig_dgrb_state.s_wait_admin~q ),
	.datab(\dgrb_state_proc~4_combout ),
	.datac(\ctrl_dgrb_r.command.cmd_tr_due~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~241_combout ),
	.cout());
defparam \sig_dgrb_state~241 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~241 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_track (
	.clk(clk),
	.d(\sig_dgrb_state~241_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_track~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_track .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_track .power_up = "low";

dffeas \sig_dgrb_last_state.s_track (
	.clk(clk),
	.d(\sig_dgrb_state.s_track~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_track~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_track .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_track .power_up = "low";

cycloneiii_lcell_comb \cdvw_proc~1 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(gnd),
	.datad(\sig_dgrb_last_state.s_track~q ),
	.cin(gnd),
	.combout(\cdvw_proc~1_combout ),
	.cout());
defparam \cdvw_proc~1 .lut_mask = 16'hEEFF;
defparam \cdvw_proc~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~430 (
	.dataa(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datab(gnd),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~430_combout ),
	.cout());
defparam \v_cdvw_state~430 .lut_mask = 16'hAFFF;
defparam \v_cdvw_state~430 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~461 (
	.dataa(\sig_cdvw_state.current_window_size[1]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~461_combout ),
	.cout());
defparam \v_cdvw_state~461 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~461 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.largest_window_size[0]~1 (
	.dataa(\sig_cdvw_state.largest_window_size[0]~0_combout ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.cout());
defparam \sig_cdvw_state.largest_window_size[0]~1 .lut_mask = 16'hFFF7;
defparam \sig_cdvw_state.largest_window_size[0]~1 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[1] (
	.clk(clk),
	.d(\v_cdvw_state~461_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[1] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[0]~6 (
	.dataa(\sig_cdvw_state.current_window_size[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~6_combout ),
	.cout(\sig_cdvw_state.current_window_size[0]~7 ));
defparam \sig_cdvw_state.current_window_size[0]~6 .lut_mask = 16'h55AA;
defparam \sig_cdvw_state.current_window_size[0]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[1]~8 (
	.dataa(\sig_cdvw_state.current_window_size[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_size[0]~7 ),
	.combout(\sig_cdvw_state.current_window_size[1]~8_combout ),
	.cout(\sig_cdvw_state.current_window_size[1]~9 ));
defparam \sig_cdvw_state.current_window_size[1]~8 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_window_size[1]~8 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \cdvw_proc~2 (
	.dataa(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector32~0_combout ),
	.cin(gnd),
	.combout(\cdvw_proc~2_combout ),
	.cout());
defparam \cdvw_proc~2 .lut_mask = 16'hAAFF;
defparam \cdvw_proc~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~530 (
	.dataa(\v_cdvw_state~529_combout ),
	.datab(\cdvw_proc~2_combout ),
	.datac(\sig_cdvw_state.working_window[63]~q ),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~530_combout ),
	.cout());
defparam \v_cdvw_state~530 .lut_mask = 16'h8BFF;
defparam \v_cdvw_state~530 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_cdvw_shift_in~4 (
	.dataa(\rsc_block:sig_chkd_all_dq_pins~q ),
	.datab(\rsc_proc~1_combout ),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\sig_rsc_cdvw_shift_in~4_combout ),
	.cout());
defparam \sig_rsc_cdvw_shift_in~4 .lut_mask = 16'hEEFF;
defparam \sig_rsc_cdvw_shift_in~4 .sum_lutc_input = "datac";

dffeas sig_rsc_cdvw_shift_in(
	.clk(clk),
	.d(\sig_rsc_cdvw_shift_in~4_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\sig_rsc_cdvw_shift_in~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_shift_in.is_wysiwyg = "true";
defparam sig_rsc_cdvw_shift_in.power_up = "low";

cycloneiii_lcell_comb \shift_in_mmc_seq_value~0 (
	.dataa(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_mmc_seq_done_1t~q ),
	.cin(gnd),
	.combout(\shift_in_mmc_seq_value~0_combout ),
	.cout());
defparam \shift_in_mmc_seq_value~0 .lut_mask = 16'hFF55;
defparam \shift_in_mmc_seq_value~0 .sum_lutc_input = "datac";

dffeas sig_trk_cdvw_shift_in(
	.clk(clk),
	.d(\shift_in_mmc_seq_value~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_shift_in~q ),
	.prn(vcc));
defparam sig_trk_cdvw_shift_in.is_wysiwyg = "true";
defparam sig_trk_cdvw_shift_in.power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.working_window[12]~4 (
	.dataa(\WideOr11~2_combout ),
	.datab(\sig_rsc_cdvw_shift_in~q ),
	.datac(\sig_dgrb_state.s_track~q ),
	.datad(\sig_trk_cdvw_shift_in~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.working_window[12]~4_combout ),
	.cout());
defparam \sig_cdvw_state.working_window[12]~4 .lut_mask = 16'hBFFF;
defparam \sig_cdvw_state.working_window[12]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.working_window[12]~5 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_cdvw_state.working_window[12]~4_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.working_window[12]~5_combout ),
	.cout());
defparam \sig_cdvw_state.working_window[12]~5 .lut_mask = 16'hAAFF;
defparam \sig_cdvw_state.working_window[12]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~531 (
	.dataa(\cdvw_proc~1_combout ),
	.datab(\v_cdvw_state~530_combout ),
	.datac(\sig_cdvw_state.working_window[12]~5_combout ),
	.datad(\sig_cdvw_state.working_window[63]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~531_combout ),
	.cout());
defparam \v_cdvw_state~531 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~531 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[63] (
	.clk(clk),
	.d(\v_cdvw_state~531_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.working_window[63]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[63] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[63] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~527 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[63]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~527_combout ),
	.cout());
defparam \v_cdvw_state~527 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~527 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.working_window[12]~6 (
	.dataa(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datab(\Selector32~0_combout ),
	.datac(\sig_cdvw_state.working_window[12]~5_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.working_window[12]~6_combout ),
	.cout());
defparam \sig_cdvw_state.working_window[12]~6 .lut_mask = 16'hFFFB;
defparam \sig_cdvw_state.working_window[12]~6 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[62] (
	.clk(clk),
	.d(\v_cdvw_state~527_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[62]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[62] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[62] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~526 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[62]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~526_combout ),
	.cout());
defparam \v_cdvw_state~526 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~526 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[61] (
	.clk(clk),
	.d(\v_cdvw_state~526_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[61]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[61] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[61] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~525 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[61]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~525_combout ),
	.cout());
defparam \v_cdvw_state~525 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~525 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[60] (
	.clk(clk),
	.d(\v_cdvw_state~525_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[60]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[60] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[60] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~524 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[60]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~524_combout ),
	.cout());
defparam \v_cdvw_state~524 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~524 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[59] (
	.clk(clk),
	.d(\v_cdvw_state~524_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[59]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[59] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[59] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~523 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[59]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~523_combout ),
	.cout());
defparam \v_cdvw_state~523 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~523 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[58] (
	.clk(clk),
	.d(\v_cdvw_state~523_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[58]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[58] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[58] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~522 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[58]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~522_combout ),
	.cout());
defparam \v_cdvw_state~522 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~522 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[57] (
	.clk(clk),
	.d(\v_cdvw_state~522_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[57]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[57] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[57] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~521 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[57]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~521_combout ),
	.cout());
defparam \v_cdvw_state~521 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~521 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[56] (
	.clk(clk),
	.d(\v_cdvw_state~521_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[56]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[56] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[56] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~520 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[56]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~520_combout ),
	.cout());
defparam \v_cdvw_state~520 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~520 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[55] (
	.clk(clk),
	.d(\v_cdvw_state~520_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[55]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[55] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[55] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~519 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[55]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~519_combout ),
	.cout());
defparam \v_cdvw_state~519 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~519 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[54] (
	.clk(clk),
	.d(\v_cdvw_state~519_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[54]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[54] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[54] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~518 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[54]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~518_combout ),
	.cout());
defparam \v_cdvw_state~518 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~518 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[53] (
	.clk(clk),
	.d(\v_cdvw_state~518_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[53]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[53] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[53] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~517 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[53]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~517_combout ),
	.cout());
defparam \v_cdvw_state~517 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~517 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[52] (
	.clk(clk),
	.d(\v_cdvw_state~517_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[52]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[52] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[52] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~516 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[52]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~516_combout ),
	.cout());
defparam \v_cdvw_state~516 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~516 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[51] (
	.clk(clk),
	.d(\v_cdvw_state~516_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[51]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[51] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[51] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~515 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[51]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~515_combout ),
	.cout());
defparam \v_cdvw_state~515 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~515 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[50] (
	.clk(clk),
	.d(\v_cdvw_state~515_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[50]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[50] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[50] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~514 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[50]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~514_combout ),
	.cout());
defparam \v_cdvw_state~514 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~514 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[49] (
	.clk(clk),
	.d(\v_cdvw_state~514_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[49]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[49] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[49] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~513 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[49]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~513_combout ),
	.cout());
defparam \v_cdvw_state~513 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~513 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[48] (
	.clk(clk),
	.d(\v_cdvw_state~513_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[48]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[48] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[48] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~512 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[48]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~512_combout ),
	.cout());
defparam \v_cdvw_state~512 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~512 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[47] (
	.clk(clk),
	.d(\v_cdvw_state~512_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[47]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[47] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[47] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~511 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[47]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~511_combout ),
	.cout());
defparam \v_cdvw_state~511 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~511 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[46] (
	.clk(clk),
	.d(\v_cdvw_state~511_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[46]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[46] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[46] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~510 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[46]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~510_combout ),
	.cout());
defparam \v_cdvw_state~510 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~510 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[45] (
	.clk(clk),
	.d(\v_cdvw_state~510_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[45]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[45] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[45] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~509 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[45]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~509_combout ),
	.cout());
defparam \v_cdvw_state~509 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~509 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[44] (
	.clk(clk),
	.d(\v_cdvw_state~509_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[44]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[44] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[44] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~508 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[44]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~508_combout ),
	.cout());
defparam \v_cdvw_state~508 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~508 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[43] (
	.clk(clk),
	.d(\v_cdvw_state~508_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[43]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[43] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[43] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~507 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[43]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~507_combout ),
	.cout());
defparam \v_cdvw_state~507 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~507 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[42] (
	.clk(clk),
	.d(\v_cdvw_state~507_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[42]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[42] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[42] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~506 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[42]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~506_combout ),
	.cout());
defparam \v_cdvw_state~506 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~506 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[41] (
	.clk(clk),
	.d(\v_cdvw_state~506_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[41]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[41] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[41] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~505 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[41]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~505_combout ),
	.cout());
defparam \v_cdvw_state~505 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~505 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[40] (
	.clk(clk),
	.d(\v_cdvw_state~505_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[40]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[40] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[40] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~504 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[40]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~504_combout ),
	.cout());
defparam \v_cdvw_state~504 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~504 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[39] (
	.clk(clk),
	.d(\v_cdvw_state~504_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[39]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[39] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[39] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~503 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[39]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~503_combout ),
	.cout());
defparam \v_cdvw_state~503 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~503 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[38] (
	.clk(clk),
	.d(\v_cdvw_state~503_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[38]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[38] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[38] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~502 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[38]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~502_combout ),
	.cout());
defparam \v_cdvw_state~502 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~502 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[37] (
	.clk(clk),
	.d(\v_cdvw_state~502_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[37]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[37] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[37] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~501 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[37]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~501_combout ),
	.cout());
defparam \v_cdvw_state~501 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~501 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[36] (
	.clk(clk),
	.d(\v_cdvw_state~501_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[36]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[36] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[36] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~500 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[36]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~500_combout ),
	.cout());
defparam \v_cdvw_state~500 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~500 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[35] (
	.clk(clk),
	.d(\v_cdvw_state~500_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[35]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[35] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[35] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~499 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[35]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~499_combout ),
	.cout());
defparam \v_cdvw_state~499 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~499 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[34] (
	.clk(clk),
	.d(\v_cdvw_state~499_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[34]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[34] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[34] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~498 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[34]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~498_combout ),
	.cout());
defparam \v_cdvw_state~498 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~498 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[33] (
	.clk(clk),
	.d(\v_cdvw_state~498_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[33]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[33] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[33] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~497 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[33]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~497_combout ),
	.cout());
defparam \v_cdvw_state~497 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~497 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[32] (
	.clk(clk),
	.d(\v_cdvw_state~497_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[32]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[32] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[32] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~496 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[32]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~496_combout ),
	.cout());
defparam \v_cdvw_state~496 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~496 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[31] (
	.clk(clk),
	.d(\v_cdvw_state~496_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[31]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[31] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[31] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~495 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[31]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~495_combout ),
	.cout());
defparam \v_cdvw_state~495 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~495 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[30] (
	.clk(clk),
	.d(\v_cdvw_state~495_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[30]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[30] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[30] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~494 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[30]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~494_combout ),
	.cout());
defparam \v_cdvw_state~494 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~494 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[29] (
	.clk(clk),
	.d(\v_cdvw_state~494_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[29]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[29] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[29] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~493 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[29]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~493_combout ),
	.cout());
defparam \v_cdvw_state~493 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~493 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[28] (
	.clk(clk),
	.d(\v_cdvw_state~493_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[28]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[28] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[28] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~492 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[28]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~492_combout ),
	.cout());
defparam \v_cdvw_state~492 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~492 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[27] (
	.clk(clk),
	.d(\v_cdvw_state~492_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[27]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[27] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[27] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~491 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[27]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~491_combout ),
	.cout());
defparam \v_cdvw_state~491 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~491 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[26] (
	.clk(clk),
	.d(\v_cdvw_state~491_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[26]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[26] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[26] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~490 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[26]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~490_combout ),
	.cout());
defparam \v_cdvw_state~490 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~490 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[25] (
	.clk(clk),
	.d(\v_cdvw_state~490_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[25]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[25] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[25] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~489 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[25]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~489_combout ),
	.cout());
defparam \v_cdvw_state~489 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~489 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[24] (
	.clk(clk),
	.d(\v_cdvw_state~489_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[24]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[24] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[24] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~488 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[24]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~488_combout ),
	.cout());
defparam \v_cdvw_state~488 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~488 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[23] (
	.clk(clk),
	.d(\v_cdvw_state~488_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[23]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[23] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[23] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~487 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[23]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~487_combout ),
	.cout());
defparam \v_cdvw_state~487 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~487 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[22] (
	.clk(clk),
	.d(\v_cdvw_state~487_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[22]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[22] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[22] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~486 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[22]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~486_combout ),
	.cout());
defparam \v_cdvw_state~486 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~486 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[21] (
	.clk(clk),
	.d(\v_cdvw_state~486_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[21]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[21] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[21] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~485 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[21]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~485_combout ),
	.cout());
defparam \v_cdvw_state~485 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~485 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[20] (
	.clk(clk),
	.d(\v_cdvw_state~485_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[20]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[20] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[20] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~484 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[20]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~484_combout ),
	.cout());
defparam \v_cdvw_state~484 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~484 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[19] (
	.clk(clk),
	.d(\v_cdvw_state~484_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[19]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[19] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[19] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~483 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[19]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~483_combout ),
	.cout());
defparam \v_cdvw_state~483 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~483 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[18] (
	.clk(clk),
	.d(\v_cdvw_state~483_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[18]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[18] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[18] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~482 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[18]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~482_combout ),
	.cout());
defparam \v_cdvw_state~482 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~482 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[17] (
	.clk(clk),
	.d(\v_cdvw_state~482_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[17]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[17] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[17] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~481 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[17]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~481_combout ),
	.cout());
defparam \v_cdvw_state~481 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~481 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[16] (
	.clk(clk),
	.d(\v_cdvw_state~481_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[16]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[16] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[16] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~480 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[16]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~480_combout ),
	.cout());
defparam \v_cdvw_state~480 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~480 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[15] (
	.clk(clk),
	.d(\v_cdvw_state~480_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[15]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[15] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[15] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~479 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[15]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~479_combout ),
	.cout());
defparam \v_cdvw_state~479 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~479 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[14] (
	.clk(clk),
	.d(\v_cdvw_state~479_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[14]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[14] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[14] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~478 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[14]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~478_combout ),
	.cout());
defparam \v_cdvw_state~478 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~478 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[13] (
	.clk(clk),
	.d(\v_cdvw_state~478_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[13]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[13] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[13] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~477 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[13]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~477_combout ),
	.cout());
defparam \v_cdvw_state~477 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~477 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[12] (
	.clk(clk),
	.d(\v_cdvw_state~477_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[12]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[12] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[12] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~476 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[12]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~476_combout ),
	.cout());
defparam \v_cdvw_state~476 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~476 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[11] (
	.clk(clk),
	.d(\v_cdvw_state~476_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[11]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[11] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[11] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~475 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[11]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~475_combout ),
	.cout());
defparam \v_cdvw_state~475 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~475 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[10] (
	.clk(clk),
	.d(\v_cdvw_state~475_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[10]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[10] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[10] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~474 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[10]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~474_combout ),
	.cout());
defparam \v_cdvw_state~474 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~474 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[9] (
	.clk(clk),
	.d(\v_cdvw_state~474_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[9]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[9] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[9] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~473 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[9]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~473_combout ),
	.cout());
defparam \v_cdvw_state~473 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~473 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[8] (
	.clk(clk),
	.d(\v_cdvw_state~473_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[8]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[8] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[8] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~472 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[8]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~472_combout ),
	.cout());
defparam \v_cdvw_state~472 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~472 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[7] (
	.clk(clk),
	.d(\v_cdvw_state~472_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[7]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[7] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[7] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~471 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[7]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~471_combout ),
	.cout());
defparam \v_cdvw_state~471 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~471 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[6] (
	.clk(clk),
	.d(\v_cdvw_state~471_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[6]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[6] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[6] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~470 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[6]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~470_combout ),
	.cout());
defparam \v_cdvw_state~470 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~470 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[5] (
	.clk(clk),
	.d(\v_cdvw_state~470_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[5] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~469 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[5]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~469_combout ),
	.cout());
defparam \v_cdvw_state~469 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~469 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[4] (
	.clk(clk),
	.d(\v_cdvw_state~469_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[4] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~468 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[4]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~468_combout ),
	.cout());
defparam \v_cdvw_state~468 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~468 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[3] (
	.clk(clk),
	.d(\v_cdvw_state~468_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[3] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~467 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[3]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~467_combout ),
	.cout());
defparam \v_cdvw_state~467 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~467 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[2] (
	.clk(clk),
	.d(\v_cdvw_state~467_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[2] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~466 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[2]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~466_combout ),
	.cout());
defparam \v_cdvw_state~466 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~466 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[1] (
	.clk(clk),
	.d(\v_cdvw_state~466_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[1] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~463 (
	.dataa(\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_dgrb_last_state.s_track~q ),
	.datad(\sig_cdvw_state.working_window[1]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~463_combout ),
	.cout());
defparam \v_cdvw_state~463 .lut_mask = 16'hFFF7;
defparam \v_cdvw_state~463 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.working_window[0] (
	.clk(clk),
	.d(\v_cdvw_state~463_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[12]~6_combout ),
	.q(\sig_cdvw_state.working_window[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[0] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~456 (
	.dataa(\sig_cdvw_state.working_window[12]~5_combout ),
	.datab(\sig_cdvw_state.last_bit_value~q ),
	.datac(\sig_cdvw_state.working_window[0]~q ),
	.datad(\v_cdvw_state~430_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~456_combout ),
	.cout());
defparam \v_cdvw_state~456 .lut_mask = 16'hFFD8;
defparam \v_cdvw_state~456 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.last_bit_value (
	.clk(clk),
	.d(\v_cdvw_state~456_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.last_bit_value~q ),
	.prn(vcc));
defparam \sig_cdvw_state.last_bit_value .is_wysiwyg = "true";
defparam \sig_cdvw_state.last_bit_value .power_up = "low";

cycloneiii_lcell_comb \find_centre_of_largest_data_valid_window~7 (
	.dataa(\sig_cdvw_state.working_window[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_cdvw_state.last_bit_value~q ),
	.cin(gnd),
	.combout(\find_centre_of_largest_data_valid_window~7_combout ),
	.cout());
defparam \find_centre_of_largest_data_valid_window~7 .lut_mask = 16'hAAFF;
defparam \find_centre_of_largest_data_valid_window~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[0]~18 (
	.dataa(\cdvw_proc~1_combout ),
	.datab(\find_centre_of_largest_data_valid_window~7_combout ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_block:sig_cdvw_calc_1t~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_size[0]~18 .lut_mask = 16'hFEFF;
defparam \sig_cdvw_state.current_window_size[0]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[0]~20 (
	.dataa(\sig_cdvw_state.current_window_size[0]~19_combout ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_size[0]~20 .lut_mask = 16'hFFF7;
defparam \sig_cdvw_state.current_window_size[0]~20 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.current_window_size[1] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[1]~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[1] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[2]~10 (
	.dataa(\sig_cdvw_state.current_window_size[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_size[1]~9 ),
	.combout(\sig_cdvw_state.current_window_size[2]~10_combout ),
	.cout(\sig_cdvw_state.current_window_size[2]~11 ));
defparam \sig_cdvw_state.current_window_size[2]~10 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_window_size[2]~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[3]~12 (
	.dataa(\sig_cdvw_state.current_window_size[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_size[2]~11 ),
	.combout(\sig_cdvw_state.current_window_size[3]~12_combout ),
	.cout(\sig_cdvw_state.current_window_size[3]~13 ));
defparam \sig_cdvw_state.current_window_size[3]~12 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_window_size[3]~12 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_window_size[3] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[3]~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[3] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~451 (
	.dataa(\sig_cdvw_state.largest_window_size[3]~q ),
	.datab(\sig_cdvw_state.largest_window_size[1]~q ),
	.datac(\sig_cdvw_state.current_window_size[1]~q ),
	.datad(\sig_cdvw_state.current_window_size[3]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~451_combout ),
	.cout());
defparam \v_cdvw_state~451 .lut_mask = 16'h6996;
defparam \v_cdvw_state~451 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~462 (
	.dataa(\sig_cdvw_state.current_window_size[0]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~462_combout ),
	.cout());
defparam \v_cdvw_state~462 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~462 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[0] (
	.clk(clk),
	.d(\v_cdvw_state~462_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[0] .power_up = "low";

dffeas \sig_cdvw_state.current_window_size[0] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[0]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[0] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[4]~14 (
	.dataa(\sig_cdvw_state.current_window_size[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_window_size[3]~13 ),
	.combout(\sig_cdvw_state.current_window_size[4]~14_combout ),
	.cout(\sig_cdvw_state.current_window_size[4]~15 ));
defparam \sig_cdvw_state.current_window_size[4]~14 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_window_size[4]~14 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_window_size[4] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[4]~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[4] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~452 (
	.dataa(\sig_cdvw_state.largest_window_size[4]~q ),
	.datab(\sig_cdvw_state.largest_window_size[0]~q ),
	.datac(\sig_cdvw_state.current_window_size[0]~q ),
	.datad(\sig_cdvw_state.current_window_size[4]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~452_combout ),
	.cout());
defparam \v_cdvw_state~452 .lut_mask = 16'h6996;
defparam \v_cdvw_state~452 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_window_size[5]~16 (
	.dataa(\sig_cdvw_state.current_window_size[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sig_cdvw_state.current_window_size[4]~15 ),
	.combout(\sig_cdvw_state.current_window_size[5]~16_combout ),
	.cout());
defparam \sig_cdvw_state.current_window_size[5]~16 .lut_mask = 16'h5A5A;
defparam \sig_cdvw_state.current_window_size[5]~16 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_window_size[5] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[5]~16_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[5] .power_up = "low";

dffeas \sig_cdvw_state.current_window_size[2] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[2]~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~18_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~20_combout ),
	.q(\sig_cdvw_state.current_window_size[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[2] .power_up = "low";

cycloneiii_lcell_comb \LessThan0~1 (
	.dataa(\sig_cdvw_state.largest_window_size[0]~q ),
	.datab(\sig_cdvw_state.current_window_size[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h00DD;
defparam \LessThan0~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~3 (
	.dataa(\sig_cdvw_state.largest_window_size[1]~q ),
	.datab(\sig_cdvw_state.current_window_size[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h00BF;
defparam \LessThan0~3 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~5 (
	.dataa(\sig_cdvw_state.largest_window_size[2]~q ),
	.datab(\sig_cdvw_state.current_window_size[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h00DF;
defparam \LessThan0~5 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~7 (
	.dataa(\sig_cdvw_state.largest_window_size[3]~q ),
	.datab(\sig_cdvw_state.current_window_size[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h00BF;
defparam \LessThan0~7 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~9 (
	.dataa(\sig_cdvw_state.largest_window_size[4]~q ),
	.datab(\sig_cdvw_state.current_window_size[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h00DF;
defparam \LessThan0~9 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \LessThan0~10 (
	.dataa(\sig_cdvw_state.largest_window_size[5]~q ),
	.datab(\sig_cdvw_state.current_window_size[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~9_cout ),
	.combout(\LessThan0~10_combout ),
	.cout());
defparam \LessThan0~10 .lut_mask = 16'hFDFD;
defparam \LessThan0~10 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \v_cdvw_state~453 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\sig_cdvw_state.working_window[0]~q ),
	.datac(\LessThan0~10_combout ),
	.datad(\sig_cdvw_state.last_bit_value~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~453_combout ),
	.cout());
defparam \v_cdvw_state~453 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~453 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~454 (
	.dataa(\v_cdvw_state~450_combout ),
	.datab(\v_cdvw_state~451_combout ),
	.datac(\v_cdvw_state~452_combout ),
	.datad(\v_cdvw_state~453_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~454_combout ),
	.cout());
defparam \v_cdvw_state~454 .lut_mask = 16'hFFFE;
defparam \v_cdvw_state~454 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~443 (
	.dataa(\sig_cdvw_state.current_bit[0]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~443_combout ),
	.cout());
defparam \v_cdvw_state~443 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~443 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \find_centre_of_largest_data_valid_window~6 (
	.dataa(\sig_cdvw_state.last_bit_value~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\find_centre_of_largest_data_valid_window~6_combout ),
	.cout());
defparam \find_centre_of_largest_data_valid_window~6 .lut_mask = 16'hAAFF;
defparam \find_centre_of_largest_data_valid_window~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~440 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.found_a_good_edge~q ),
	.datac(\sig_cdvw_state.status.calculating~q ),
	.datad(\find_centre_of_largest_data_valid_window~6_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~440_combout ),
	.cout());
defparam \v_cdvw_state~440 .lut_mask = 16'hFFFE;
defparam \v_cdvw_state~440 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.found_a_good_edge (
	.clk(clk),
	.d(\v_cdvw_state~440_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.found_a_good_edge~q ),
	.prn(vcc));
defparam \sig_cdvw_state.found_a_good_edge .is_wysiwyg = "true";
defparam \sig_cdvw_state.found_a_good_edge .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.first_good_edge[1]~0 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.found_a_good_edge~q ),
	.datac(\sig_cdvw_state.status.calculating~q ),
	.datad(\find_centre_of_largest_data_valid_window~6_combout ),
	.cin(gnd),
	.combout(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.cout());
defparam \sig_cdvw_state.first_good_edge[1]~0 .lut_mask = 16'hFFF7;
defparam \sig_cdvw_state.first_good_edge[1]~0 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_good_edge[0] (
	.clk(clk),
	.d(\v_cdvw_state~443_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[0] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[1]~11 (
	.dataa(\sig_cdvw_state.current_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_bit[0]~7 ),
	.combout(\sig_cdvw_state.current_bit[1]~11_combout ),
	.cout(\sig_cdvw_state.current_bit[1]~12 ));
defparam \sig_cdvw_state.current_bit[1]~11 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_bit[1]~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[2]~13 (
	.dataa(\sig_cdvw_state.current_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_bit[1]~12 ),
	.combout(\sig_cdvw_state.current_bit[2]~13_combout ),
	.cout(\sig_cdvw_state.current_bit[2]~14 ));
defparam \sig_cdvw_state.current_bit[2]~13 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_bit[2]~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[5]~10 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\cdvw_proc~1_combout ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_block:sig_cdvw_calc_1t~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~10_combout ),
	.cout());
defparam \sig_cdvw_state.current_bit[5]~10 .lut_mask = 16'hFEFF;
defparam \sig_cdvw_state.current_bit[5]~10 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.current_bit[2] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[2]~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[2] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[3]~15 (
	.dataa(\sig_cdvw_state.current_bit[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_bit[2]~14 ),
	.combout(\sig_cdvw_state.current_bit[3]~15_combout ),
	.cout(\sig_cdvw_state.current_bit[3]~16 ));
defparam \sig_cdvw_state.current_bit[3]~15 .lut_mask = 16'h5A5F;
defparam \sig_cdvw_state.current_bit[3]~15 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_bit[3] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[3]~15_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[3] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[5]~8 (
	.dataa(\sig_cdvw_state.current_bit[0]~q ),
	.datab(\sig_cdvw_state.current_bit[1]~q ),
	.datac(\sig_cdvw_state.current_bit[2]~q ),
	.datad(\sig_cdvw_state.current_bit[3]~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~8_combout ),
	.cout());
defparam \sig_cdvw_state.current_bit[5]~8 .lut_mask = 16'h7FFF;
defparam \sig_cdvw_state.current_bit[5]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[4]~17 (
	.dataa(\sig_cdvw_state.current_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sig_cdvw_state.current_bit[3]~16 ),
	.combout(\sig_cdvw_state.current_bit[4]~17_combout ),
	.cout(\sig_cdvw_state.current_bit[4]~18 ));
defparam \sig_cdvw_state.current_bit[4]~17 .lut_mask = 16'h5AAF;
defparam \sig_cdvw_state.current_bit[4]~17 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_bit[4] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[4]~17_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[4] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[5]~19 (
	.dataa(\sig_cdvw_state.current_bit[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sig_cdvw_state.current_bit[4]~18 ),
	.combout(\sig_cdvw_state.current_bit[5]~19_combout ),
	.cout());
defparam \sig_cdvw_state.current_bit[5]~19 .lut_mask = 16'h5A5A;
defparam \sig_cdvw_state.current_bit[5]~19 .sum_lutc_input = "cin";

dffeas \sig_cdvw_state.current_bit[5] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[5]~19_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[5] .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.current_bit[5]~9 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.current_bit[5]~8_combout ),
	.datac(\sig_cdvw_state.current_bit[4]~q ),
	.datad(\sig_cdvw_state.current_bit[5]~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~9_combout ),
	.cout());
defparam \sig_cdvw_state.current_bit[5]~9 .lut_mask = 16'hFFF7;
defparam \sig_cdvw_state.current_bit[5]~9 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.current_bit[1] (
	.clk(clk),
	.d(\sig_cdvw_state.current_bit[1]~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~9_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~10_combout ),
	.q(\sig_cdvw_state.current_bit[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[1] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~444 (
	.dataa(\sig_cdvw_state.current_bit[1]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~444_combout ),
	.cout());
defparam \v_cdvw_state~444 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~444 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_good_edge[1] (
	.clk(clk),
	.d(\v_cdvw_state~444_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[1] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~425 (
	.dataa(\sig_cdvw_state.current_bit[0]~q ),
	.datab(\sig_cdvw_state.first_good_edge[0]~q ),
	.datac(\sig_cdvw_state.current_bit[1]~q ),
	.datad(\sig_cdvw_state.first_good_edge[1]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~425_combout ),
	.cout());
defparam \v_cdvw_state~425 .lut_mask = 16'h6996;
defparam \v_cdvw_state~425 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~445 (
	.dataa(\sig_cdvw_state.current_bit[3]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~445_combout ),
	.cout());
defparam \v_cdvw_state~445 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~445 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_good_edge[3] (
	.clk(clk),
	.d(\v_cdvw_state~445_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[3] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~446 (
	.dataa(\sig_cdvw_state.current_bit[4]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~446_combout ),
	.cout());
defparam \v_cdvw_state~446 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~446 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_good_edge[4] (
	.clk(clk),
	.d(\v_cdvw_state~446_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[1]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[4] .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~426 (
	.dataa(\sig_cdvw_state.current_bit[3]~q ),
	.datab(\sig_cdvw_state.first_good_edge[3]~q ),
	.datac(\sig_cdvw_state.current_bit[4]~q ),
	.datad(\sig_cdvw_state.first_good_edge[4]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~426_combout ),
	.cout());
defparam \v_cdvw_state~426 .lut_mask = 16'h6996;
defparam \v_cdvw_state~426 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~427 (
	.dataa(\v_cdvw_state~424_combout ),
	.datab(\v_cdvw_state~425_combout ),
	.datac(\v_cdvw_state~426_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\v_cdvw_state~427_combout ),
	.cout());
defparam \v_cdvw_state~427 .lut_mask = 16'hFEFE;
defparam \v_cdvw_state~427 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~448 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\sig_cdvw_state.valid_phase_seen~q ),
	.datac(\sig_cdvw_state.status.calculating~q ),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~448_combout ),
	.cout());
defparam \v_cdvw_state~448 .lut_mask = 16'hFEFF;
defparam \v_cdvw_state~448 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.valid_phase_seen (
	.clk(clk),
	.d(\v_cdvw_state~448_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.valid_phase_seen~q ),
	.prn(vcc));
defparam \sig_cdvw_state.valid_phase_seen .is_wysiwyg = "true";
defparam \sig_cdvw_state.valid_phase_seen .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~428 (
	.dataa(\sig_cdvw_state.invalid_phase_seen~q ),
	.datab(\sig_cdvw_state.valid_phase_seen~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\v_cdvw_state~428_combout ),
	.cout());
defparam \v_cdvw_state~428 .lut_mask = 16'hEEEE;
defparam \v_cdvw_state~428 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~449 (
	.dataa(\sig_cdvw_state.first_cycle~q ),
	.datab(\sig_cdvw_state.status.calculating~q ),
	.datac(\cdvw_proc~2_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~449_combout ),
	.cout());
defparam \v_cdvw_state~449 .lut_mask = 16'hBFFF;
defparam \v_cdvw_state~449 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.first_cycle (
	.clk(clk),
	.d(\v_cdvw_state~449_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.first_cycle~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_cycle .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_cycle .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~429 (
	.dataa(\find_centre_of_largest_data_valid_window~0_combout ),
	.datab(\v_cdvw_state~427_combout ),
	.datac(\v_cdvw_state~428_combout ),
	.datad(\sig_cdvw_state.first_cycle~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~429_combout ),
	.cout());
defparam \v_cdvw_state~429 .lut_mask = 16'h27FF;
defparam \v_cdvw_state~429 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~433 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\v_cdvw_state~429_combout ),
	.datac(\cdvw_proc~2_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~433_combout ),
	.cout());
defparam \v_cdvw_state~433 .lut_mask = 16'hBFFF;
defparam \v_cdvw_state~433 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.status.calculating (
	.clk(clk),
	.d(\v_cdvw_state~433_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.calculating~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.calculating .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.calculating .power_up = "low";

cycloneiii_lcell_comb \sig_cdvw_state.largest_window_size[0]~0 (
	.dataa(\sig_cdvw_state.last_bit_value~q ),
	.datab(\sig_cdvw_state.status.calculating~q ),
	.datac(\LessThan0~10_combout ),
	.datad(\sig_cdvw_state.working_window[0]~q ),
	.cin(gnd),
	.combout(\sig_cdvw_state.largest_window_size[0]~0_combout ),
	.cout());
defparam \sig_cdvw_state.largest_window_size[0]~0 .lut_mask = 16'hBFFF;
defparam \sig_cdvw_state.largest_window_size[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~455 (
	.dataa(\v_cdvw_state~430_combout ),
	.datab(\v_cdvw_state~454_combout ),
	.datac(\sig_cdvw_state.multiple_eq_windows~q ),
	.datad(\sig_cdvw_state.largest_window_size[0]~0_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~455_combout ),
	.cout());
defparam \v_cdvw_state~455 .lut_mask = 16'hFFFE;
defparam \v_cdvw_state~455 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.multiple_eq_windows (
	.clk(clk),
	.d(\v_cdvw_state~455_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.multiple_eq_windows~q ),
	.prn(vcc));
defparam \sig_cdvw_state.multiple_eq_windows .is_wysiwyg = "true";
defparam \sig_cdvw_state.multiple_eq_windows .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~431 (
	.dataa(\find_centre_of_largest_data_valid_window~0_combout ),
	.datab(\sig_cdvw_state.multiple_eq_windows~q ),
	.datac(\sig_cdvw_state.status.valid_result~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\v_cdvw_state~431_combout ),
	.cout());
defparam \v_cdvw_state~431 .lut_mask = 16'hFF96;
defparam \v_cdvw_state~431 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~432 (
	.dataa(\v_cdvw_state~429_combout ),
	.datab(\v_cdvw_state~430_combout ),
	.datac(\sig_cdvw_state.status.valid_result~q ),
	.datad(\v_cdvw_state~431_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~432_combout ),
	.cout());
defparam \v_cdvw_state~432 .lut_mask = 16'hEDDE;
defparam \v_cdvw_state~432 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.status.valid_result (
	.clk(clk),
	.d(\v_cdvw_state~432_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.valid_result~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.valid_result .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.valid_result .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~127 (
	.dataa(\Selector127~1_combout ),
	.datab(\sig_cdvw_state.status.valid_result~q ),
	.datac(seq_ac_add_1t_ac_lat_internal),
	.datad(\sig_dgrb_state.s_track~q ),
	.cin(gnd),
	.combout(\sig_trk_state~127_combout ),
	.cout());
defparam \sig_trk_state~127 .lut_mask = 16'hBFFF;
defparam \sig_trk_state~127 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_idle (
	.clk(clk),
	.d(\sig_trk_state~127_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_idle~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_idle .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_idle .power_up = "low";

cycloneiii_lcell_comb \Selector123~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector123~0_combout ),
	.cout());
defparam \Selector123~0 .lut_mask = 16'hAAFF;
defparam \Selector123~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector86~0 (
	.dataa(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(\shift_in_mmc_seq_value~0_combout ),
	.datac(\Equal10~0_combout ),
	.datad(\Equal10~1_combout ),
	.cin(gnd),
	.combout(\Selector86~0_combout ),
	.cout());
defparam \Selector86~0 .lut_mask = 16'hBFFF;
defparam \Selector86~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~128 (
	.dataa(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(\Equal10~0_combout ),
	.datac(\Equal10~1_combout ),
	.datad(\shift_in_mmc_seq_value~0_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~128_combout ),
	.cout());
defparam \sig_trk_state~128 .lut_mask = 16'hFFBF;
defparam \sig_trk_state~128 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~121 (
	.dataa(\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_state~121_combout ),
	.cout());
defparam \sig_trk_state~121 .lut_mask = 16'hEEEE;
defparam \sig_trk_state~121 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~122 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_state~121_combout ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(\sig_trk_state~113_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~122_combout ),
	.cout());
defparam \sig_trk_state~122 .lut_mask = 16'hFFFE;
defparam \sig_trk_state~122 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_wait (
	.clk(clk),
	.d(\sig_trk_state~122_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_wait .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_wait .power_up = "low";

cycloneiii_lcell_comb \sig_phs_shft_end~0 (
	.dataa(\sig_phs_shft_busy~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.cin(gnd),
	.combout(\sig_phs_shft_end~0_combout ),
	.cout());
defparam \sig_phs_shft_end~0 .lut_mask = 16'hAAFF;
defparam \sig_phs_shft_end~0 .sum_lutc_input = "datac";

dffeas sig_phs_shft_end(
	.clk(clk),
	.d(\sig_phs_shft_end~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_end~q ),
	.prn(vcc));
defparam sig_phs_shft_end.is_wysiwyg = "true";
defparam sig_phs_shft_end.power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~109 (
	.dataa(\sig_cdvw_state.status.calculating~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datad(\sig_phs_shft_end~q ),
	.cin(gnd),
	.combout(\sig_trk_state~109_combout ),
	.cout());
defparam \sig_trk_state~109 .lut_mask = 16'h8BFF;
defparam \sig_trk_state~109 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_last_state~29 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_last_state~29_combout ),
	.cout());
defparam \sig_trk_last_state~29 .lut_mask = 16'hEEEE;
defparam \sig_trk_last_state~29 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_last_state.s_trk_cdvw_drift (
	.clk(clk),
	.d(\sig_trk_last_state~29_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_drift .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_drift .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~107 (
	.dataa(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datab(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_state~107_combout ),
	.cout());
defparam \sig_trk_state~107 .lut_mask = 16'hEEEE;
defparam \sig_trk_state~107 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~114 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_state~107_combout ),
	.datac(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(\sig_trk_state~113_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~114_combout ),
	.cout());
defparam \sig_trk_state~114 .lut_mask = 16'hFFFE;
defparam \sig_trk_state~114 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_adjust_resync (
	.clk(clk),
	.d(\sig_trk_state~114_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_adjust_resync .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_adjust_resync .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~108 (
	.dataa(\sig_trk_state~106_combout ),
	.datab(gnd),
	.datac(\sig_phs_shft_end~q ),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\sig_trk_state~108_combout ),
	.cout());
defparam \sig_trk_state~108 .lut_mask = 16'hAFFF;
defparam \sig_trk_state~108 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_last_state~30 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_last_state~30_combout ),
	.cout());
defparam \sig_trk_last_state~30 .lut_mask = 16'hEEEE;
defparam \sig_trk_last_state~30 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_last_state.s_trk_cdvw_calc (
	.clk(clk),
	.d(\sig_trk_last_state~30_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_calc .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_calc .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~110 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\sig_trk_state~110_combout ),
	.cout());
defparam \sig_trk_state~110 .lut_mask = 16'hBFFF;
defparam \sig_trk_state~110 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~117 (
	.dataa(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datab(\sig_phs_shft_end~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datad(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.cin(gnd),
	.combout(\sig_trk_state~117_combout ),
	.cout());
defparam \sig_trk_state~117 .lut_mask = 16'h53FF;
defparam \sig_trk_state~117 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~118 (
	.dataa(\Selector86~0_combout ),
	.datab(\sig_trk_state~117_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.cin(gnd),
	.combout(\sig_trk_state~118_combout ),
	.cout());
defparam \sig_trk_state~118 .lut_mask = 16'hEEFF;
defparam \sig_trk_state~118 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector127~1 (
	.dataa(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\Selector127~1_combout ),
	.cout());
defparam \Selector127~1 .lut_mask = 16'hAAFF;
defparam \Selector127~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~119 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\sig_trk_state~110_combout ),
	.datac(\sig_trk_state~118_combout ),
	.datad(\Selector127~1_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~119_combout ),
	.cout());
defparam \sig_trk_state~119 .lut_mask = 16'hFAFC;
defparam \sig_trk_state~119 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector93~0 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector93~0_combout ),
	.cout());
defparam \Selector93~0 .lut_mask = 16'hEEEE;
defparam \Selector93~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_mimic_cdv[0]~0 (
	.dataa(\sig_cdvw_state.status.valid_result~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\trk_block:sig_mimic_cdv[0]~0_combout ),
	.cout());
defparam \trk_block:sig_mimic_cdv[0]~0 .lut_mask = 16'hEEEE;
defparam \trk_block:sig_mimic_cdv[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector93~1 (
	.dataa(\trk_block:sig_mimic_cdv_found~q ),
	.datab(\Selector93~0_combout ),
	.datac(\trk_block:sig_mimic_cdv[0]~0_combout ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\Selector93~1_combout ),
	.cout());
defparam \Selector93~1 .lut_mask = 16'hFEFF;
defparam \Selector93~1 .sum_lutc_input = "datac";

dffeas \trk_block:sig_mimic_cdv_found (
	.clk(clk),
	.d(\Selector93~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_mimic_cdv_found~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv_found .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv_found .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~123 (
	.dataa(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datab(\trk_block:sig_mimic_cdv_found~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\sig_trk_state~123_combout ),
	.cout());
defparam \sig_trk_state~123 .lut_mask = 16'hEFFE;
defparam \sig_trk_state~123 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~124 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_state~108_combout ),
	.datac(\sig_trk_state~119_combout ),
	.datad(\sig_trk_state~123_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~124_combout ),
	.cout());
defparam \sig_trk_state~124 .lut_mask = 16'hFFFE;
defparam \sig_trk_state~124 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_drift (
	.clk(clk),
	.d(\sig_trk_state~124_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_drift .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_drift .power_up = "low";

cycloneiii_lcell_comb \sig_trk_state~111 (
	.dataa(\sig_trk_state~110_combout ),
	.datab(gnd),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datad(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.cin(gnd),
	.combout(\sig_trk_state~111_combout ),
	.cout());
defparam \sig_trk_state~111 .lut_mask = 16'hAFFF;
defparam \sig_trk_state~111 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~112 (
	.dataa(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(\Equal10~0_combout ),
	.datac(\Equal10~1_combout ),
	.datad(\shift_in_mmc_seq_value~0_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~112_combout ),
	.cout());
defparam \sig_trk_state~112 .lut_mask = 16'hFFFE;
defparam \sig_trk_state~112 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~113 (
	.dataa(\sig_trk_state~108_combout ),
	.datab(\sig_trk_state~109_combout ),
	.datac(\sig_trk_state~111_combout ),
	.datad(\sig_trk_state~112_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~113_combout ),
	.cout());
defparam \sig_trk_state~113 .lut_mask = 16'hFEFF;
defparam \sig_trk_state~113 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~115 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_state~128_combout ),
	.datac(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datad(\sig_trk_state~113_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~115_combout ),
	.cout());
defparam \sig_trk_state~115 .lut_mask = 16'hFFFE;
defparam \sig_trk_state~115 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_next_phase (
	.clk(clk),
	.d(\sig_trk_state~115_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_next_phase .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_next_phase .power_up = "low";

cycloneiii_lcell_comb \Selector86~1 (
	.dataa(\trk_block:sig_trk_state.s_trk_idle~q ),
	.datab(\Selector86~0_combout ),
	.datac(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datad(\sig_phs_shft_end~q ),
	.cin(gnd),
	.combout(\Selector86~1_combout ),
	.cout());
defparam \Selector86~1 .lut_mask = 16'hFFFE;
defparam \Selector86~1 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_mimic_sample (
	.clk(clk),
	.d(\Selector86~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_mimic_sample .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_mimic_sample .power_up = "low";

dffeas \trk_block:trk_proc:v_remaining_samples[2] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[2]~0_combout ),
	.asdata(\Selector123~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[2]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[2] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[2] .power_up = "low";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[1]~0 (
	.dataa(\Add10~2_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[1]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[1]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[1]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[1]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector124~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector124~0_combout ),
	.cout());
defparam \Selector124~0 .lut_mask = 16'hAAFF;
defparam \Selector124~0 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[1] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[1]~0_combout ),
	.asdata(\Selector124~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[1]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[1] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[1] .power_up = "low";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[0]~0 (
	.dataa(\Add10~0_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[0]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[0]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[0]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector125~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector125~0_combout ),
	.cout());
defparam \Selector125~0 .lut_mask = 16'hAAFF;
defparam \Selector125~0 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[0] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[0]~0_combout ),
	.asdata(\Selector125~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[0]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[0] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[0] .power_up = "low";

cycloneiii_lcell_comb \Equal10~1 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[3]~q ),
	.datab(\trk_block:trk_proc:v_remaining_samples[2]~q ),
	.datac(\trk_block:trk_proc:v_remaining_samples[1]~q ),
	.datad(\trk_block:trk_proc:v_remaining_samples[0]~q ),
	.cin(gnd),
	.combout(\Equal10~1_combout ),
	.cout());
defparam \Equal10~1 .lut_mask = 16'h7FFF;
defparam \Equal10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_remaining_samples~18 (
	.dataa(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.datab(\trk_block:sig_mmc_seq_done_1t~q ),
	.datac(\Equal10~0_combout ),
	.datad(\Equal10~1_combout ),
	.cin(gnd),
	.combout(\v_remaining_samples~18_combout ),
	.cout());
defparam \v_remaining_samples~18 .lut_mask = 16'hFFFB;
defparam \v_remaining_samples~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[7]~0 (
	.dataa(\Add10~14_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[7]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[7]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[7]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[7]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector118~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector118~0_combout ),
	.cout());
defparam \Selector118~0 .lut_mask = 16'hAAFF;
defparam \Selector118~0 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[7] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[7]~0_combout ),
	.asdata(\Selector118~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[7]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[7] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[7] .power_up = "low";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[5]~0 (
	.dataa(\Add10~10_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[5]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[5]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[5]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[5]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector120~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector120~0_combout ),
	.cout());
defparam \Selector120~0 .lut_mask = 16'hAAFF;
defparam \Selector120~0 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[5] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[5]~0_combout ),
	.asdata(\Selector120~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[5]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[5] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[5] .power_up = "low";

cycloneiii_lcell_comb \trk_block:trk_proc:v_remaining_samples[4]~0 (
	.dataa(\Add10~8_combout ),
	.datab(\trk_block:trk_proc:v_remaining_samples[4]~q ),
	.datac(gnd),
	.datad(\v_remaining_samples~18_combout ),
	.cin(gnd),
	.combout(\trk_block:trk_proc:v_remaining_samples[4]~0_combout ),
	.cout());
defparam \trk_block:trk_proc:v_remaining_samples[4]~0 .lut_mask = 16'hAACC;
defparam \trk_block:trk_proc:v_remaining_samples[4]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector121~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_idle~q ),
	.cin(gnd),
	.combout(\Selector121~0_combout ),
	.cout());
defparam \Selector121~0 .lut_mask = 16'hAAFF;
defparam \Selector121~0 .sum_lutc_input = "datac";

dffeas \trk_block:trk_proc:v_remaining_samples[4] (
	.clk(clk),
	.d(\trk_block:trk_proc:v_remaining_samples[4]~0_combout ),
	.asdata(\Selector121~0_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:trk_proc:v_remaining_samples[4]~q ),
	.prn(vcc));
defparam \trk_block:trk_proc:v_remaining_samples[4] .is_wysiwyg = "true";
defparam \trk_block:trk_proc:v_remaining_samples[4] .power_up = "low";

cycloneiii_lcell_comb \Equal10~0 (
	.dataa(\trk_block:trk_proc:v_remaining_samples[6]~q ),
	.datab(\trk_block:trk_proc:v_remaining_samples[7]~q ),
	.datac(\trk_block:trk_proc:v_remaining_samples[5]~q ),
	.datad(\trk_block:trk_proc:v_remaining_samples[4]~q ),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
defparam \Equal10~0 .lut_mask = 16'h7FFF;
defparam \Equal10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~125 (
	.dataa(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(\Equal10~0_combout ),
	.datac(\Equal10~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_state~125_combout ),
	.cout());
defparam \sig_trk_state~125 .lut_mask = 16'hFEFE;
defparam \sig_trk_state~125 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~126 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datac(\sig_trk_state~125_combout ),
	.datad(\sig_trk_state~113_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~126_combout ),
	.cout());
defparam \sig_trk_state~126 .lut_mask = 16'hFAFC;
defparam \sig_trk_state~126 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_calc (
	.clk(clk),
	.d(\sig_trk_state~126_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_calc .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_calc .power_up = "low";

cycloneiii_lcell_comb \sig_trk_cdvw_calc~4 (
	.dataa(\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.cin(gnd),
	.combout(\sig_trk_cdvw_calc~4_combout ),
	.cout());
defparam \sig_trk_cdvw_calc~4 .lut_mask = 16'hFF55;
defparam \sig_trk_cdvw_calc~4 .sum_lutc_input = "datac";

dffeas sig_trk_cdvw_calc(
	.clk(clk),
	.d(\sig_trk_cdvw_calc~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_calc~q ),
	.prn(vcc));
defparam sig_trk_cdvw_calc.is_wysiwyg = "true";
defparam sig_trk_cdvw_calc.power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~258 (
	.dataa(last_states_rrp_seek),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~258_combout ),
	.cout());
defparam \sig_dgrb_state~258 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~258 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_seek_cdvw (
	.clk(clk),
	.d(\sig_dgrb_state~258_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_seek_cdvw~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_seek_cdvw .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_seek_cdvw .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~274 (
	.dataa(last_states_read_mtp),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~274_combout ),
	.cout());
defparam \sig_dgrb_state~274 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~274 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_read_mtp (
	.clk(clk),
	.d(\sig_dgrb_state~274_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_read_mtp~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_read_mtp .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_read_mtp .power_up = "low";

cycloneiii_lcell_comb \sig_rsc_req~29 (
	.dataa(\sig_rsc_ack~q ),
	.datab(gnd),
	.datac(\sig_dgrb_state.s_seek_cdvw~q ),
	.datad(\sig_dgrb_state.s_read_mtp~q ),
	.cin(gnd),
	.combout(\sig_rsc_req~29_combout ),
	.cout());
defparam \sig_rsc_req~29 .lut_mask = 16'hFFF5;
defparam \sig_rsc_req~29 .sum_lutc_input = "datac";

dffeas \sig_rsc_req.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\sig_rsc_req~29_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_cdvw_calc .power_up = "low";

cycloneiii_lcell_comb \Selector55~0 (
	.dataa(\Selector49~0_combout ),
	.datab(\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.datad(\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.cin(gnd),
	.combout(\Selector55~0_combout ),
	.cout());
defparam \Selector55~0 .lut_mask = 16'hFEFF;
defparam \Selector55~0 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\Selector55~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_calc .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc .power_up = "low";

cycloneiii_lcell_comb \Selector55~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.cin(gnd),
	.combout(\Selector55~1_combout ),
	.cout());
defparam \Selector55~1 .lut_mask = 16'hAAFF;
defparam \Selector55~1 .sum_lutc_input = "datac";

dffeas sig_rsc_cdvw_calc(
	.clk(clk),
	.d(\Selector55~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_calc.is_wysiwyg = "true";
defparam sig_rsc_cdvw_calc.power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~260 (
	.dataa(last_states_rrp_sweep),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~260_combout ),
	.cout());
defparam \sig_dgrb_state~260 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~260 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_test_phases (
	.clk(clk),
	.d(\sig_dgrb_state~260_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_test_phases~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_test_phases .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_test_phases .power_up = "low";

cycloneiii_lcell_comb \WideOr11~2 (
	.dataa(gnd),
	.datab(\sig_dgrb_state.s_seek_cdvw~q ),
	.datac(\sig_dgrb_state.s_test_phases~q ),
	.datad(\sig_dgrb_state.s_read_mtp~q ),
	.cin(gnd),
	.combout(\WideOr11~2_combout ),
	.cout());
defparam \WideOr11~2 .lut_mask = 16'h3FFF;
defparam \WideOr11~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector32~0 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_trk_cdvw_calc~q ),
	.datac(\sig_rsc_cdvw_calc~q ),
	.datad(\WideOr11~2_combout ),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'hFEFF;
defparam \Selector32~0 .sum_lutc_input = "datac";

dffeas \cdvw_block:sig_cdvw_calc_1t (
	.clk(clk),
	.d(\Selector32~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cdvw_block:sig_cdvw_calc_1t~q ),
	.prn(vcc));
defparam \cdvw_block:sig_cdvw_calc_1t .is_wysiwyg = "true";
defparam \cdvw_block:sig_cdvw_calc_1t .power_up = "low";

cycloneiii_lcell_comb \v_cdvw_state~439 (
	.dataa(\sig_cdvw_state.current_window_centre[0]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~439_combout ),
	.cout());
defparam \v_cdvw_state~439 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~439 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_centre[0] (
	.clk(clk),
	.d(\v_cdvw_state~439_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_centre[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[0] .power_up = "low";

cycloneiii_lcell_comb \Selector74~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\sig_cdvw_state.largest_window_centre[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector74~0_combout ),
	.cout());
defparam \Selector74~0 .lut_mask = 16'hEEEE;
defparam \Selector74~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~1 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~1_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~1 .lut_mask = 16'hAAFF;
defparam \rsc_block:sig_count[6]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[5]~1 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[5]~1_combout ),
	.cout());
defparam \rsc_block:sig_count[5]~1 .lut_mask = 16'hEFFF;
defparam \rsc_block:sig_count[5]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[5]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datad(\rsc_block:sig_count[5]~1_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[5]~2_combout ),
	.cout());
defparam \rsc_block:sig_count[5]~2 .lut_mask = 16'h0FFF;
defparam \rsc_block:sig_count[5]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector46~0 (
	.dataa(\sig_cdvw_state.largest_window_centre[0]~q ),
	.datab(\Add6~0_combout ),
	.datac(\rsc_block:sig_count[6]~1_combout ),
	.datad(\rsc_block:sig_count[5]~2_combout ),
	.cin(gnd),
	.combout(\Selector46~0_combout ),
	.cout());
defparam \Selector46~0 .lut_mask = 16'hACFF;
defparam \Selector46~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[6]~5 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsc_block:sig_count[6]~5_combout ),
	.cout());
defparam \rsc_block:sig_count[6]~5 .lut_mask = 16'hEEEE;
defparam \rsc_block:sig_count[6]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[5]~3 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsc_block:sig_count[5]~3_combout ),
	.cout());
defparam \rsc_block:sig_count[5]~3 .lut_mask = 16'hEEEE;
defparam \rsc_block:sig_count[5]~3 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw .power_up = "low";

cycloneiii_lcell_comb \Selector69~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector69~0_combout ),
	.cout());
defparam \Selector69~0 .lut_mask = 16'hEEEE;
defparam \Selector69~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \WideOr13~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\WideOr13~1_combout ),
	.cout());
defparam \WideOr13~1 .lut_mask = 16'hBFFF;
defparam \WideOr13~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[5]~0 (
	.dataa(\sig_phs_shft_end~q ),
	.datab(\Equal7~2_combout ),
	.datac(\Selector69~0_combout ),
	.datad(\WideOr13~1_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[5]~0_combout ),
	.cout());
defparam \rsc_block:sig_count[5]~0 .lut_mask = 16'hBFFF;
defparam \rsc_block:sig_count[5]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \rsc_block:sig_count[5]~4 (
	.dataa(\rsc_block:sig_count[6]~3_combout ),
	.datab(\rsc_block:sig_count[6]~5_combout ),
	.datac(\rsc_block:sig_count[5]~3_combout ),
	.datad(\rsc_block:sig_count[5]~0_combout ),
	.cin(gnd),
	.combout(\rsc_block:sig_count[5]~4_combout ),
	.cout());
defparam \rsc_block:sig_count[5]~4 .lut_mask = 16'hFF7F;
defparam \rsc_block:sig_count[5]~4 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_count[0] (
	.clk(clk),
	.d(\Selector46~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[5]~4_combout ),
	.q(\rsc_block:sig_count[0]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[0] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[0] .power_up = "low";

cycloneiii_lcell_comb \Equal7~2 (
	.dataa(\Equal7~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\rsc_block:sig_count[0]~q ),
	.cin(gnd),
	.combout(\Equal7~2_combout ),
	.cout());
defparam \Equal7~2 .lut_mask = 16'hAAFF;
defparam \Equal7~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector57~1 (
	.dataa(\Selector57~0_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(\Equal7~2_combout ),
	.datad(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.cin(gnd),
	.combout(\Selector57~1_combout ),
	.cout());
defparam \Selector57~1 .lut_mask = 16'hEFFF;
defparam \Selector57~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_seek_cdvw (
	.clk(clk),
	.d(\Selector57~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_seek_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_seek_cdvw .power_up = "low";

cycloneiii_lcell_comb \Selector69~3 (
	.dataa(\Selector69~1_combout ),
	.datab(\sig_cdvw_state.status.valid_result~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.cin(gnd),
	.combout(\Selector69~3_combout ),
	.cout());
defparam \Selector69~3 .lut_mask = 16'hFEFF;
defparam \Selector69~3 .sum_lutc_input = "datac";

dffeas \cal_codvw_phase[0] (
	.clk(clk),
	.d(\Selector74~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector69~3_combout ),
	.q(\cal_codvw_phase[0]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[0] .is_wysiwyg = "true";
defparam \cal_codvw_phase[0] .power_up = "low";

cycloneiii_lcell_comb \Add5~8 (
	.dataa(\Add5~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_num_phase_shifts[0]~q ),
	.datad(\Add9~0_combout ),
	.cin(gnd),
	.combout(\Add5~8_combout ),
	.cout());
defparam \Add5~8 .lut_mask = 16'h8BFF;
defparam \Add5~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add5~11 (
	.dataa(\Add5~7_combout ),
	.datab(\Add5~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~10 ),
	.combout(\Add5~11_combout ),
	.cout(\Add5~12 ));
defparam \Add5~11 .lut_mask = 16'h96DF;
defparam \Add5~11 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add5~25 (
	.dataa(\Add9~2_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~11_combout ),
	.cin(gnd),
	.combout(\Add5~25_combout ),
	.cout());
defparam \Add5~25 .lut_mask = 16'h47FF;
defparam \Add5~25 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_num_phase_shifts[1] (
	.clk(clk),
	.d(\Add5~25_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[1]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[1] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[1] .power_up = "low";

cycloneiii_lcell_comb \Equal6~1 (
	.dataa(\Equal6~0_combout ),
	.datab(gnd),
	.datac(\rsc_block:sig_num_phase_shifts[1]~q ),
	.datad(\rsc_block:sig_num_phase_shifts[0]~q ),
	.cin(gnd),
	.combout(\Equal6~1_combout ),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hAFFF;
defparam \Equal6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~0 (
	.dataa(\rsc_block:sig_chkd_all_dq_pins~q ),
	.datab(\Selector51~0_combout ),
	.datac(gnd),
	.datad(\Equal6~1_combout ),
	.cin(gnd),
	.combout(\Selector53~0_combout ),
	.cout());
defparam \Selector53~0 .lut_mask = 16'hEEFF;
defparam \Selector53~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector53~1 (
	.dataa(\Selector59~0_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Selector53~0_combout ),
	.cin(gnd),
	.combout(\Selector53~1_combout ),
	.cout());
defparam \Selector53~1 .lut_mask = 16'hFFFE;
defparam \Selector53~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_rewind_phase (
	.clk(clk),
	.d(\Selector53~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_rewind_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_rewind_phase .power_up = "low";

cycloneiii_lcell_comb \Selector69~1 (
	.dataa(\Equal7~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datad(\rsc_block:sig_count[0]~q ),
	.cin(gnd),
	.combout(\Selector69~1_combout ),
	.cout());
defparam \Selector69~1 .lut_mask = 16'hFEFF;
defparam \Selector69~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector83~4 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datab(\sig_dgrb_state.s_read_mtp~q ),
	.datac(\sig_cdvw_state.status.valid_result~q ),
	.datad(\sig_cdvw_state.status.calculating~q ),
	.cin(gnd),
	.combout(\Selector83~4_combout ),
	.cout());
defparam \Selector83~4 .lut_mask = 16'hEFFF;
defparam \Selector83~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector83~5 (
	.dataa(\Equal6~1_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(\Selector69~1_combout ),
	.datad(\Selector83~4_combout ),
	.cin(gnd),
	.combout(\Selector83~5_combout ),
	.cout());
defparam \Selector83~5 .lut_mask = 16'hFFFD;
defparam \Selector83~5 .sum_lutc_input = "datac";

dffeas sig_rsc_ack(
	.clk(clk),
	.d(\Selector83~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_ack~q ),
	.prn(vcc));
defparam sig_rsc_ack.is_wysiwyg = "true";
defparam sig_rsc_ack.power_up = "low";

cycloneiii_lcell_comb \Selector23~0 (
	.dataa(\sig_dgrb_state.s_test_phases~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_rsc_ack~q ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
defparam \Selector23~0 .lut_mask = 16'hAAFF;
defparam \Selector23~0 .sum_lutc_input = "datac";

dffeas \sig_rsc_req.s_rsc_test_phase (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_test_phase~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_test_phase .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_test_phase .power_up = "low";

cycloneiii_lcell_comb \Selector47~0 (
	.dataa(gnd),
	.datab(\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.datac(\sig_rsc_req.s_rsc_test_phase~q ),
	.datad(\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.cin(gnd),
	.combout(\Selector47~0_combout ),
	.cout());
defparam \Selector47~0 .lut_mask = 16'h3FFF;
defparam \Selector47~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector47~1 (
	.dataa(\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.datab(\Selector47~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datad(\Selector83~5_combout ),
	.cin(gnd),
	.combout(\Selector47~1_combout ),
	.cout());
defparam \Selector47~1 .lut_mask = 16'hF7FF;
defparam \Selector47~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_idle (
	.clk(clk),
	.d(\Selector47~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_idle .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_idle .power_up = "low";

cycloneiii_lcell_comb \Selector49~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datad(\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.cin(gnd),
	.combout(\Selector49~0_combout ),
	.cout());
defparam \Selector49~0 .lut_mask = 16'h0FFF;
defparam \Selector49~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector49~1 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datab(\Selector49~0_combout ),
	.datac(\sig_rsc_req.s_rsc_test_phase~q ),
	.datad(\sig_phs_shft_end~q ),
	.cin(gnd),
	.combout(\Selector49~1_combout ),
	.cout());
defparam \Selector49~1 .lut_mask = 16'hFFFE;
defparam \Selector49~1 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_test_phase (
	.clk(clk),
	.d(\Selector49~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_test_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_test_phase .power_up = "low";

dffeas \ctrl_dgrb_r.command_op.single_bit (
	.clk(clk),
	.d(\ctrl_dgrb.command_op.single_bit ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command_op.single_bit~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command_op.single_bit .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command_op.single_bit .power_up = "low";

dffeas single_bit_cal(
	.clk(clk),
	.d(\ctrl_dgrb_r.command_op.single_bit~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ac_muxctrl_broadcast_rcommand_req),
	.q(\single_bit_cal~q ),
	.prn(vcc));
defparam single_bit_cal.is_wysiwyg = "true";
defparam single_bit_cal.power_up = "low";

cycloneiii_lcell_comb \Selector38~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datac(\sig_dq_pin_ctr[0]~q ),
	.datad(\single_bit_cal~q ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hEFFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

dffeas \sig_dq_pin_ctr[0] (
	.clk(clk),
	.d(\Selector38~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dq_pin_ctr[3]~16_combout ),
	.q(\sig_dq_pin_ctr[0]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[0] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[0] .power_up = "low";

cycloneiii_lcell_comb \Mux1~2 (
	.dataa(\sig_dq_pin_ctr[3]~q ),
	.datab(q_b_14),
	.datac(\sig_dq_pin_ctr[2]~q ),
	.datad(q_b_10),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hFFDE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~3 (
	.dataa(q_b_26),
	.datab(\sig_dq_pin_ctr[3]~q ),
	.datac(\Mux1~2_combout ),
	.datad(q_b_30),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hFFBE;
defparam \Mux1~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~4 (
	.dataa(\sig_dq_pin_ctr[2]~q ),
	.datab(q_b_24),
	.datac(\sig_dq_pin_ctr[3]~q ),
	.datad(q_b_8),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'hFFDE;
defparam \Mux1~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~5 (
	.dataa(q_b_12),
	.datab(\sig_dq_pin_ctr[2]~q ),
	.datac(\Mux1~4_combout ),
	.datad(q_b_28),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hFFBE;
defparam \Mux1~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~6 (
	.dataa(\sig_dq_pin_ctr[0]~q ),
	.datab(\Mux1~3_combout ),
	.datac(\sig_dq_pin_ctr[1]~q ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
defparam \Mux1~6 .lut_mask = 16'hFFDE;
defparam \Mux1~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~7 (
	.dataa(\sig_dq_pin_ctr[3]~q ),
	.datab(q_b_15),
	.datac(\sig_dq_pin_ctr[2]~q ),
	.datad(q_b_11),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
defparam \Mux1~7 .lut_mask = 16'hFFDE;
defparam \Mux1~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~8 (
	.dataa(q_b_27),
	.datab(\sig_dq_pin_ctr[3]~q ),
	.datac(\Mux1~7_combout ),
	.datad(q_b_31),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
defparam \Mux1~8 .lut_mask = 16'hFFBE;
defparam \Mux1~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Mux1~9 (
	.dataa(\Mux1~1_combout ),
	.datab(\sig_dq_pin_ctr[0]~q ),
	.datac(\Mux1~6_combout ),
	.datad(\Mux1~8_combout ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
defparam \Mux1~9 .lut_mask = 16'hFFBE;
defparam \Mux1~9 .sum_lutc_input = "datac";

dffeas \tp_match_block:sig_rdata_current_pin[15] (
	.clk(clk),
	.d(\Mux1~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[15] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[15] .power_up = "low";

cycloneiii_lcell_comb \Equal9~0 (
	.dataa(\Equal8~0_combout ),
	.datab(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.datac(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal9~0_combout ),
	.cout());
defparam \Equal9~0 .lut_mask = 16'hFEFE;
defparam \Equal9~0 .sum_lutc_input = "datac";

dffeas sig_poa_match(
	.clk(clk),
	.d(\Equal9~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_match~q ),
	.prn(vcc));
defparam sig_poa_match.is_wysiwyg = "true";
defparam sig_poa_match.power_up = "low";

dffeas \tp_match_block:sig_rdata_valid_1t (
	.clk(clk),
	.d(rdata_valid[0]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_valid_1t~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_valid_1t .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_valid_1t .power_up = "low";

cycloneiii_lcell_comb \poa_match_proc~0 (
	.dataa(\tp_match_block:sig_rdata_valid_2t~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\tp_match_block:sig_rdata_valid_1t~q ),
	.cin(gnd),
	.combout(\poa_match_proc~0_combout ),
	.cout());
defparam \poa_match_proc~0 .lut_mask = 16'hAAFF;
defparam \poa_match_proc~0 .sum_lutc_input = "datac";

dffeas sig_poa_match_en(
	.clk(clk),
	.d(\poa_match_proc~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_match_en~q ),
	.prn(vcc));
defparam sig_poa_match_en.is_wysiwyg = "true";
defparam sig_poa_match_en.power_up = "low";

cycloneiii_lcell_comb \sig_poa_state~4 (
	.dataa(\sig_dgrb_state.s_poa_cal~q ),
	.datab(\poa_block:sig_poa_state~q ),
	.datac(\sig_poa_match~q ),
	.datad(\sig_poa_match_en~q ),
	.cin(gnd),
	.combout(\sig_poa_state~4_combout ),
	.cout());
defparam \sig_poa_state~4 .lut_mask = 16'hFFFE;
defparam \sig_poa_state~4 .sum_lutc_input = "datac";

dffeas \poa_block:sig_poa_state (
	.clk(clk),
	.d(\sig_poa_state~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\poa_block:sig_poa_state~q ),
	.prn(vcc));
defparam \poa_block:sig_poa_state .is_wysiwyg = "true";
defparam \poa_block:sig_poa_state .power_up = "low";

cycloneiii_lcell_comb \sig_poa_ack~3 (
	.dataa(\sig_dgrb_state.s_poa_cal~q ),
	.datab(\poa_block:sig_poa_state~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_poa_ack~3_combout ),
	.cout());
defparam \sig_poa_ack~3 .lut_mask = 16'hEEEE;
defparam \sig_poa_ack~3 .sum_lutc_input = "datac";

dffeas sig_poa_ack(
	.clk(clk),
	.d(\sig_poa_ack~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_ack~q ),
	.prn(vcc));
defparam sig_poa_ack.is_wysiwyg = "true";
defparam sig_poa_ack.power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~246 (
	.dataa(\sig_trk_ack~q ),
	.datab(\sig_poa_ack~q ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_track~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~246_combout ),
	.cout());
defparam \sig_dgrb_state~246 .lut_mask = 16'hAACC;
defparam \sig_dgrb_state~246 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~247 (
	.dataa(\sig_dgrb_state~245_combout ),
	.datab(\sig_dgrb_state~246_combout ),
	.datac(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datad(\sig_dgrb_state.s_adv_rd_lat~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~247_combout ),
	.cout());
defparam \sig_dgrb_state~247 .lut_mask = 16'hEFFF;
defparam \sig_dgrb_state~247 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_req~27 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sig_dgrb_state.s_seek_cdvw~q ),
	.datad(\sig_dgrb_state.s_read_mtp~q ),
	.cin(gnd),
	.combout(\sig_rsc_req~27_combout ),
	.cout());
defparam \sig_rsc_req~27 .lut_mask = 16'h0FFF;
defparam \sig_rsc_req~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~242 (
	.dataa(\sig_rsc_ack~q ),
	.datab(\sig_dgrb_state.s_reset_cdvw~q ),
	.datac(\sig_dgrb_state.s_test_phases~q ),
	.datad(\sig_rsc_req~27_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~242_combout ),
	.cout());
defparam \sig_dgrb_state~242 .lut_mask = 16'hFEFF;
defparam \sig_dgrb_state~242 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~270 (
	.dataa(\sig_dgrb_state.s_release_admin~q ),
	.datab(\sig_dgrb_state~247_combout ),
	.datac(\sig_dgrb_state~261_combout ),
	.datad(\sig_dgrb_state~242_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~270_combout ),
	.cout());
defparam \sig_dgrb_state~270 .lut_mask = 16'h27FF;
defparam \sig_dgrb_state~270 .sum_lutc_input = "datac";

dffeas \sig_dgrb_last_state.s_adv_wd_lat (
	.clk(clk),
	.d(\sig_dgrb_state.s_adv_wd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_adv_wd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_adv_wd_lat .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~251 (
	.dataa(\sig_dgrb_state~249_combout ),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~251_combout ),
	.cout());
defparam \sig_dgrb_state~251 .lut_mask = 16'hACFF;
defparam \sig_dgrb_state~251 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~255 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datad(\sig_dgrb_state.s_wait_admin~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~255_combout ),
	.cout());
defparam \sig_dgrb_state~255 .lut_mask = 16'h0FFF;
defparam \sig_dgrb_state~255 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~271 (
	.dataa(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(\sig_dgrb_state~251_combout ),
	.datad(\sig_dgrb_state~255_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~271_combout ),
	.cout());
defparam \sig_dgrb_state~271 .lut_mask = 16'hBFFF;
defparam \sig_dgrb_state~271 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~272 (
	.dataa(\sig_dgrb_state~266_combout ),
	.datab(\sig_dgrb_state~269_combout ),
	.datac(\sig_dgrb_state~270_combout ),
	.datad(\sig_dgrb_state~271_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~272_combout ),
	.cout());
defparam \sig_dgrb_state~272 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~272 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_adv_rd_lat (
	.clk(clk),
	.d(\sig_dgrb_state~272_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_adv_rd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_rd_lat .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~254 (
	.dataa(\sig_dgrb_state~253_combout ),
	.datab(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datac(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datad(\sig_dgrb_state.s_adv_rd_lat~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~254_combout ),
	.cout());
defparam \sig_dgrb_state~254 .lut_mask = 16'hBFFF;
defparam \sig_dgrb_state~254 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~256 (
	.dataa(\sig_dgrb_state~255_combout ),
	.datab(ac_muxctrl_broadcast_rcommand_req),
	.datac(\sig_dgrb_state.s_idle~q ),
	.datad(\sig_dgrb_state.s_release_admin~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~256_combout ),
	.cout());
defparam \sig_dgrb_state~256 .lut_mask = 16'hFEFF;
defparam \sig_dgrb_state~256 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~257 (
	.dataa(\sig_dgrb_state~250_combout ),
	.datab(\sig_dgrb_state~254_combout ),
	.datac(\sig_dgrb_state~256_combout ),
	.datad(\sig_dgrb_state.s_wait_admin~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~257_combout ),
	.cout());
defparam \sig_dgrb_state~257 .lut_mask = 16'h7FFF;
defparam \sig_dgrb_state~257 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~263 (
	.dataa(\dgrb_state_proc~4_combout ),
	.datab(\sig_dgrb_state~262_combout ),
	.datac(\sig_dgrb_state~257_combout ),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~263_combout ),
	.cout());
defparam \sig_dgrb_state~263 .lut_mask = 16'hFF7F;
defparam \sig_dgrb_state~263 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_idle (
	.clk(clk),
	.d(\sig_dgrb_state~263_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_idle .power_up = "low";

cycloneiii_lcell_comb \dgrb_state_proc~4 (
	.dataa(curr_cmdcmd_idle),
	.datab(\sig_dgrb_state.s_release_admin~q ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\dgrb_state_proc~4_combout ),
	.cout());
defparam \dgrb_state_proc~4 .lut_mask = 16'hEEFF;
defparam \dgrb_state_proc~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~265 (
	.dataa(last_states_adv_rd_lat),
	.datab(\sig_dgrb_state.s_wait_admin~q ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_dgrb_state~265_combout ),
	.cout());
defparam \sig_dgrb_state~265 .lut_mask = 16'hFEFE;
defparam \sig_dgrb_state~265 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_adv_rd_lat_setup (
	.clk(clk),
	.d(\sig_dgrb_state~265_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state~281_combout ),
	.q(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_rd_lat_setup .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_rd_lat_setup .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~243 (
	.dataa(sig_doing_rd_0),
	.datab(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~243_combout ),
	.cout());
defparam \sig_dgrb_state~243 .lut_mask = 16'hEEFF;
defparam \sig_dgrb_state~243 .sum_lutc_input = "datac";

dffeas \sig_dgrb_last_state.s_adv_rd_lat_setup (
	.clk(clk),
	.d(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_adv_rd_lat_setup .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_adv_rd_lat_setup .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~267 (
	.dataa(\dgrb_state_proc~4_combout ),
	.datab(gnd),
	.datac(\sig_dgrb_state~243_combout ),
	.datad(\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~267_combout ),
	.cout());
defparam \sig_dgrb_state~267 .lut_mask = 16'hAFFF;
defparam \sig_dgrb_state~267 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~239 (
	.dataa(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~239_combout ),
	.cout());
defparam \sig_dgrb_state~239 .lut_mask = 16'hAAFF;
defparam \sig_dgrb_state~239 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~273 (
	.dataa(\sig_dgrb_state~268_combout ),
	.datab(\sig_dgrb_state~267_combout ),
	.datac(\sig_dgrb_state.s_wait_admin~q ),
	.datad(\sig_dgrb_state~239_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~273_combout ),
	.cout());
defparam \sig_dgrb_state~273 .lut_mask = 16'hEFFF;
defparam \sig_dgrb_state~273 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_wait_admin (
	.clk(clk),
	.d(\sig_dgrb_state~273_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_wait_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_wait_admin .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_wait_admin .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~238 (
	.dataa(last_states_rdv),
	.datab(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_wait_admin~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~238_combout ),
	.cout());
defparam \sig_dgrb_state~238 .lut_mask = 16'hAACC;
defparam \sig_dgrb_state~238 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~240 (
	.dataa(\dgrb_state_proc~4_combout ),
	.datab(\sig_dgrb_state~237_combout ),
	.datac(\sig_dgrb_state~238_combout ),
	.datad(\sig_dgrb_state~239_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~240_combout ),
	.cout());
defparam \sig_dgrb_state~240 .lut_mask = 16'hFAFC;
defparam \sig_dgrb_state~240 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_rdata_valid_align (
	.clk(clk),
	.d(\sig_dgrb_state~240_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_rdata_valid_align~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_rdata_valid_align .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_rdata_valid_align .power_up = "low";

cycloneiii_lcell_comb \sig_dgrb_state~277 (
	.dataa(\sig_dgrb_state.s_adv_rd_lat~q ),
	.datab(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datac(q_b_0),
	.datad(q_b_8),
	.cin(gnd),
	.combout(\sig_dgrb_state~277_combout ),
	.cout());
defparam \sig_dgrb_state~277 .lut_mask = 16'hEFFF;
defparam \sig_dgrb_state~277 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~278 (
	.dataa(\seq_rdata_valid_lat_dec~3_combout ),
	.datab(\sig_dgrb_state~277_combout ),
	.datac(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datad(\sig_dgrb_state.s_adv_wd_lat~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~278_combout ),
	.cout());
defparam \sig_dgrb_state~278 .lut_mask = 16'hFFFE;
defparam \sig_dgrb_state~278 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~282 (
	.dataa(\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(\sig_dgrb_state.s_read_mtp~q ),
	.datac(\sig_dgrb_state.s_reset_cdvw~q ),
	.datad(\sig_dgrb_state.s_test_phases~q ),
	.cin(gnd),
	.combout(\sig_dgrb_state~282_combout ),
	.cout());
defparam \sig_dgrb_state~282 .lut_mask = 16'h7FFF;
defparam \sig_dgrb_state~282 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~279 (
	.dataa(\sig_rsc_ack~q ),
	.datab(\sig_dgrb_state.s_release_admin~q ),
	.datac(\sig_dgrb_state~261_combout ),
	.datad(\sig_dgrb_state~282_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~279_combout ),
	.cout());
defparam \sig_dgrb_state~279 .lut_mask = 16'hEFFF;
defparam \sig_dgrb_state~279 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_dgrb_state~280 (
	.dataa(\sig_dgrb_state~276_combout ),
	.datab(\sig_dgrb_state~278_combout ),
	.datac(\dgrb_state_proc~4_combout ),
	.datad(\sig_dgrb_state~279_combout ),
	.cin(gnd),
	.combout(\sig_dgrb_state~280_combout ),
	.cout());
defparam \sig_dgrb_state~280 .lut_mask = 16'hFFEF;
defparam \sig_dgrb_state~280 .sum_lutc_input = "datac";

dffeas \sig_dgrb_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgrb_state~280_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_release_admin .power_up = "low";

cycloneiii_lcell_comb \Selector21~1 (
	.dataa(\Selector21~0_combout ),
	.datab(\sig_dgrb_state.s_release_admin~q ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
defparam \Selector21~1 .lut_mask = 16'hFF77;
defparam \Selector21~1 .sum_lutc_input = "datac";

dffeas \sig_ac_req.s_ac_idle (
	.clk(clk),
	.d(\Selector21~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_idle~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_idle .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_idle .power_up = "low";

cycloneiii_lcell_comb \Selector24~0 (
	.dataa(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datab(\sig_dgrb_state.s_adv_rd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hEEEE;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector25~1 (
	.dataa(\Selector25~0_combout ),
	.datab(\sig_dgrb_state.s_test_phases~q ),
	.datac(\sig_rsc_ack~q ),
	.datad(\sig_rsc_req~27_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
defparam \Selector25~1 .lut_mask = 16'hFEFF;
defparam \Selector25~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector24~1 (
	.dataa(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(\Selector24~0_combout ),
	.datac(\sig_ac_req.s_ac_read_rdv~q ),
	.datad(\Selector25~1_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
defparam \Selector24~1 .lut_mask = 16'hFFFE;
defparam \Selector24~1 .sum_lutc_input = "datac";

dffeas \sig_ac_req.s_ac_read_rdv (
	.clk(clk),
	.d(\Selector24~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_rdv .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_rdv .power_up = "low";

cycloneiii_lcell_comb \sig_addr_cmd_state~39 (
	.dataa(\sig_addr_cmd_state~38_combout ),
	.datab(\sig_ac_req.s_ac_read_rdv~q ),
	.datac(\WideOr26~2_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~39_combout ),
	.cout());
defparam \sig_addr_cmd_state~39 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd_state~39 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_rdv (
	.clk(clk),
	.d(\sig_addr_cmd_state~39_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_rdv .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_rdv .power_up = "low";

cycloneiii_lcell_comb \WideOr26~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(\sig_ac_req.s_ac_read_rdv~q ),
	.datad(\sig_ac_req.s_ac_read_mtp~q ),
	.cin(gnd),
	.combout(\WideOr26~1_combout ),
	.cout());
defparam \WideOr26~1 .lut_mask = 16'h6996;
defparam \WideOr26~1 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv .power_up = "low";

cycloneiii_lcell_comb \Selector175~10 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector175~10_combout ),
	.cout());
defparam \Selector175~10 .lut_mask = 16'hEEEE;
defparam \Selector175~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector25~2 (
	.dataa(\sig_dgrb_state.s_poa_cal~q ),
	.datab(\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datac(\Selector25~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
defparam \Selector25~2 .lut_mask = 16'hFEFE;
defparam \Selector25~2 .sum_lutc_input = "datac";

dffeas \sig_ac_req.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\Selector25~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_poa_mtp .power_up = "low";

cycloneiii_lcell_comb \sig_addr_cmd_state~42 (
	.dataa(\sig_addr_cmd_state~38_combout ),
	.datab(\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datac(\WideOr26~2_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~42_combout ),
	.cout());
defparam \sig_addr_cmd_state~42 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd_state~42 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\sig_addr_cmd_state~42_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp .power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_relax (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_relax .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_relax .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_count[7]~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~1_combout ),
	.cout());
defparam \ac_block:sig_count[7]~1 .lut_mask = 16'hAAFF;
defparam \ac_block:sig_count[7]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[7]~2 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(\Equal13~1_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datad(\ac_block:sig_count[7]~1_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~2_combout ),
	.cout());
defparam \ac_block:sig_count[7]~2 .lut_mask = 16'hBFFF;
defparam \ac_block:sig_count[7]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[5]~2 (
	.dataa(\ac_block:sig_count[5]~1_combout ),
	.datab(\Equal13~1_combout ),
	.datac(\Selector175~10_combout ),
	.datad(\ac_block:sig_count[7]~2_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[5]~2_combout ),
	.cout());
defparam \ac_block:sig_count[5]~2 .lut_mask = 16'hFEFF;
defparam \ac_block:sig_count[5]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector168~0 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(\Equal13~1_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(\ac_block:sig_count[7]~1_combout ),
	.cin(gnd),
	.combout(\Selector168~0_combout ),
	.cout());
defparam \Selector168~0 .lut_mask = 16'hBFFF;
defparam \Selector168~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[7]~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~0_combout ),
	.cout());
defparam \ac_block:sig_count[7]~0 .lut_mask = 16'hAAFF;
defparam \ac_block:sig_count[7]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector173~0 (
	.dataa(\Add23~0_combout ),
	.datab(\ac_block:sig_count[5]~2_combout ),
	.datac(\Selector168~0_combout ),
	.datad(\ac_block:sig_count[7]~0_combout ),
	.cin(gnd),
	.combout(\Selector173~0_combout ),
	.cout());
defparam \Selector173~0 .lut_mask = 16'h8BFF;
defparam \Selector173~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[5]~0 (
	.dataa(\ac_block:sig_count[7]~6_combout ),
	.datab(\Equal13~1_combout ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[5]~0_combout ),
	.cout());
defparam \ac_block:sig_count[5]~0 .lut_mask = 16'hFEFF;
defparam \ac_block:sig_count[5]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[5]~3 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[5]~3_combout ),
	.cout());
defparam \ac_block:sig_count[5]~3 .lut_mask = 16'h6996;
defparam \ac_block:sig_count[5]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[5]~4 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_count[5]~0_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(\ac_block:sig_count[5]~3_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[5]~4_combout ),
	.cout());
defparam \ac_block:sig_count[5]~4 .lut_mask = 16'h7FF7;
defparam \ac_block:sig_count[5]~4 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[0] (
	.clk(clk),
	.d(\Selector173~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[5]~4_combout ),
	.q(\ac_block:sig_count[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[0] .is_wysiwyg = "true";
defparam \ac_block:sig_count[0] .power_up = "low";

cycloneiii_lcell_comb \sig_burst_count~4 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\sig_burst_count~4_combout ),
	.cout());
defparam \sig_burst_count~4 .lut_mask = 16'hFF77;
defparam \sig_burst_count~4 .sum_lutc_input = "datac";

dffeas \ac_block:sig_burst_count[0] (
	.clk(clk),
	.d(\sig_burst_count~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_burst_count[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_burst_count[0] .is_wysiwyg = "true";
defparam \ac_block:sig_burst_count[0] .power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_count[7]~4 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~4_combout ),
	.cout());
defparam \ac_block:sig_count[7]~4 .lut_mask = 16'hAACC;
defparam \ac_block:sig_count[7]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[1]~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac_block:sig_count[1]~0_combout ),
	.cout());
defparam \ac_block:sig_count[1]~0 .lut_mask = 16'hEEEE;
defparam \ac_block:sig_count[1]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[7]~7 (
	.dataa(\ac_block:sig_count[5]~0_combout ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(\ac_block:sig_count[7]~4_combout ),
	.datad(\ac_block:sig_count[1]~0_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~7_combout ),
	.cout());
defparam \ac_block:sig_count[7]~7 .lut_mask = 16'hFF7F;
defparam \ac_block:sig_count[7]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[1]~1 (
	.dataa(\ac_block:sig_count[7]~1_combout ),
	.datab(\ac_block:sig_count[1]~0_combout ),
	.datac(\Equal13~1_combout ),
	.datad(\ac_block:sig_count[7]~4_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[1]~1_combout ),
	.cout());
defparam \ac_block:sig_count[1]~1 .lut_mask = 16'hFEFF;
defparam \ac_block:sig_count[1]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[1]~2 (
	.dataa(\Add23~2_combout ),
	.datab(\ac_block:sig_count[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac_block:sig_count[1]~2_combout ),
	.cout());
defparam \ac_block:sig_count[1]~2 .lut_mask = 16'hEEEE;
defparam \ac_block:sig_count[1]~2 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_count[7]~8 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(\Equal13~1_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~8_combout ),
	.cout());
defparam \ac_block:sig_count[7]~8 .lut_mask = 16'hEEFF;
defparam \ac_block:sig_count[7]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_count[1]~3 (
	.dataa(\ac_block:sig_count[1]~q ),
	.datab(\ac_block:sig_count[7]~7_combout ),
	.datac(\ac_block:sig_count[1]~2_combout ),
	.datad(\ac_block:sig_count[7]~8_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[1]~3_combout ),
	.cout());
defparam \ac_block:sig_count[1]~3 .lut_mask = 16'hB8FF;
defparam \ac_block:sig_count[1]~3 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[1] (
	.clk(clk),
	.d(\ac_block:sig_count[1]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_count[1]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[1] .is_wysiwyg = "true";
defparam \ac_block:sig_count[1] .power_up = "low";

cycloneiii_lcell_comb \Equal13~1 (
	.dataa(\Equal13~0_combout ),
	.datab(gnd),
	.datac(\ac_block:sig_count[0]~q ),
	.datad(\ac_block:sig_count[1]~q ),
	.cin(gnd),
	.combout(\Equal13~1_combout ),
	.cout());
defparam \Equal13~1 .lut_mask = 16'hAFFF;
defparam \Equal13~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd_state~38 (
	.dataa(gnd),
	.datab(\Equal13~1_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~38_combout ),
	.cout());
defparam \sig_addr_cmd_state~38 .lut_mask = 16'h3FFF;
defparam \sig_addr_cmd_state~38 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd_state~44 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datab(\sig_addr_cmd_state~38_combout ),
	.datac(gnd),
	.datad(\WideOr26~2_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~44_combout ),
	.cout());
defparam \sig_addr_cmd_state~44 .lut_mask = 16'hEEFF;
defparam \sig_addr_cmd_state~44 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_relax (
	.clk(clk),
	.d(\sig_addr_cmd_state~44_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_relax .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_relax .power_up = "low";

cycloneiii_lcell_comb \WideOr26~2 (
	.dataa(\WideOr26~0_combout ),
	.datab(\WideOr26~1_combout ),
	.datac(\sig_ac_req.s_ac_idle~q ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\WideOr26~2_combout ),
	.cout());
defparam \WideOr26~2 .lut_mask = 16'hFEFF;
defparam \WideOr26~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd_state~43 (
	.dataa(\sig_addr_cmd_state~38_combout ),
	.datab(\sig_ac_req.s_ac_idle~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datad(\WideOr26~2_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~43_combout ),
	.cout());
defparam \sig_addr_cmd_state~43 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd_state~43 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_idle (
	.clk(clk),
	.d(\sig_addr_cmd_state~43_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_idle .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_idle .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_setup[0]~1 (
	.dataa(\ac_block:sig_setup[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac_block:sig_setup[0]~1_combout ),
	.cout(\ac_block:sig_setup[0]~2 ));
defparam \ac_block:sig_setup[0]~1 .lut_mask = 16'h5555;
defparam \ac_block:sig_setup[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_setup[1]~1 (
	.dataa(\ac_block:sig_setup[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_block:sig_setup[0]~2 ),
	.combout(\ac_block:sig_setup[1]~1_combout ),
	.cout(\ac_block:sig_setup[1]~2 ));
defparam \ac_block:sig_setup[1]~1 .lut_mask = 16'h5AAF;
defparam \ac_block:sig_setup[1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \ac_block:sig_setup[2]~1 (
	.dataa(\ac_block:sig_setup[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_block:sig_setup[1]~2 ),
	.combout(\ac_block:sig_setup[2]~1_combout ),
	.cout(\ac_block:sig_setup[2]~2 ));
defparam \ac_block:sig_setup[2]~1 .lut_mask = 16'h5A5F;
defparam \ac_block:sig_setup[2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \ac_block:sig_setup[3]~1 (
	.dataa(\ac_block:sig_setup[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_block:sig_setup[2]~2 ),
	.combout(\ac_block:sig_setup[3]~1_combout ),
	.cout(\ac_block:sig_setup[3]~2 ));
defparam \ac_block:sig_setup[3]~1 .lut_mask = 16'h5AAF;
defparam \ac_block:sig_setup[3]~1 .sum_lutc_input = "cin";

dffeas \ac_block:sig_setup[3] (
	.clk(clk),
	.d(\ac_block:sig_setup[3]~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!dgb_ac_access_gnt_r),
	.ena(\ac_block:sig_setup[4]~1_combout ),
	.q(\ac_block:sig_setup[3]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[3] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[3] .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_setup[4]~2 (
	.dataa(\ac_block:sig_setup[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ac_block:sig_setup[3]~2 ),
	.combout(\ac_block:sig_setup[4]~2_combout ),
	.cout());
defparam \ac_block:sig_setup[4]~2 .lut_mask = 16'h5A5A;
defparam \ac_block:sig_setup[4]~2 .sum_lutc_input = "cin";

dffeas \ac_block:sig_setup[4] (
	.clk(clk),
	.d(\ac_block:sig_setup[4]~2_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!dgb_ac_access_gnt_r),
	.ena(\ac_block:sig_setup[4]~1_combout ),
	.q(\ac_block:sig_setup[4]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[4] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[4] .power_up = "low";

cycloneiii_lcell_comb \dimm_driving_dq_proc~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\dimm_driving_dq_proc~1_combout ),
	.cout());
defparam \dimm_driving_dq_proc~1 .lut_mask = 16'hAAFF;
defparam \dimm_driving_dq_proc~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_block:sig_setup[4]~1 (
	.dataa(\Selector128~0_combout ),
	.datab(\ac_block:sig_setup[3]~q ),
	.datac(\ac_block:sig_setup[4]~q ),
	.datad(\dimm_driving_dq_proc~1_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_setup[4]~1_combout ),
	.cout());
defparam \ac_block:sig_setup[4]~1 .lut_mask = 16'hFF7F;
defparam \ac_block:sig_setup[4]~1 .sum_lutc_input = "datac";

dffeas \ac_block:sig_setup[0] (
	.clk(clk),
	.d(\ac_block:sig_setup[0]~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!dgb_ac_access_gnt_r),
	.ena(\ac_block:sig_setup[4]~1_combout ),
	.q(\ac_block:sig_setup[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[0] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[0] .power_up = "low";

dffeas \ac_block:sig_setup[1] (
	.clk(clk),
	.d(\ac_block:sig_setup[1]~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!dgb_ac_access_gnt_r),
	.ena(\ac_block:sig_setup[4]~1_combout ),
	.q(\ac_block:sig_setup[1]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[1] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[1] .power_up = "low";

dffeas \ac_block:sig_setup[2] (
	.clk(clk),
	.d(\ac_block:sig_setup[2]~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!dgb_ac_access_gnt_r),
	.ena(\ac_block:sig_setup[4]~1_combout ),
	.q(\ac_block:sig_setup[2]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[2] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[2] .power_up = "low";

cycloneiii_lcell_comb \Selector128~0 (
	.dataa(dgb_ac_access_gnt_r),
	.datab(\ac_block:sig_setup[0]~q ),
	.datac(\ac_block:sig_setup[1]~q ),
	.datad(\ac_block:sig_setup[2]~q ),
	.cin(gnd),
	.combout(\Selector128~0_combout ),
	.cout());
defparam \Selector128~0 .lut_mask = 16'hFFFE;
defparam \Selector128~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector128~1 (
	.dataa(\ac_block:sig_setup[3]~q ),
	.datab(\ac_block:sig_setup[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector128~1_combout ),
	.cout());
defparam \Selector128~1 .lut_mask = 16'hEEEE;
defparam \Selector128~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector128~2 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datac(\Selector128~0_combout ),
	.datad(\Selector128~1_combout ),
	.cin(gnd),
	.combout(\Selector128~2_combout ),
	.cout());
defparam \Selector128~2 .lut_mask = 16'h7FFF;
defparam \Selector128~2 .sum_lutc_input = "datac";

dffeas sig_dimm_driving_dq(
	.clk(clk),
	.d(\Selector128~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dimm_driving_dq~q ),
	.prn(vcc));
defparam sig_dimm_driving_dq.is_wysiwyg = "true";
defparam sig_dimm_driving_dq.power_up = "low";

cycloneiii_lcell_comb \Selector52~0 (
	.dataa(\Equal7~1_combout ),
	.datab(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datac(\sig_dimm_driving_dq~q ),
	.datad(\rsc_block:sig_count[0]~q ),
	.cin(gnd),
	.combout(\Selector52~0_combout ),
	.cout());
defparam \Selector52~0 .lut_mask = 16'hEFFF;
defparam \Selector52~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector51~3 (
	.dataa(\Selector51~2_combout ),
	.datab(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datac(gnd),
	.datad(\Selector52~0_combout ),
	.cin(gnd),
	.combout(\Selector51~3_combout ),
	.cout());
defparam \Selector51~3 .lut_mask = 16'hEEFF;
defparam \Selector51~3 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_rsc_state.s_rsc_flush_datapath (
	.clk(clk),
	.d(\Selector51~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_flush_datapath .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_flush_datapath .power_up = "low";

cycloneiii_lcell_comb \WideOr13~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.cin(gnd),
	.combout(\WideOr13~0_combout ),
	.cout());
defparam \WideOr13~0 .lut_mask = 16'hFFF0;
defparam \WideOr13~0 .sum_lutc_input = "datac";

dffeas sig_rsc_ac_access_req(
	.clk(clk),
	.d(\WideOr13~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_ac_access_req~q ),
	.prn(vcc));
defparam sig_rsc_ac_access_req.is_wysiwyg = "true";
defparam sig_rsc_ac_access_req.power_up = "low";

cycloneiii_lcell_comb \Selector23~1 (
	.dataa(\sig_ac_req.s_ac_read_mtp~q ),
	.datab(\sig_rsc_ac_access_req~q ),
	.datac(\Selector23~0_combout ),
	.datad(\Selector25~1_combout ),
	.cin(gnd),
	.combout(\Selector23~1_combout ),
	.cout());
defparam \Selector23~1 .lut_mask = 16'hFFFE;
defparam \Selector23~1 .sum_lutc_input = "datac";

dffeas \sig_ac_req.s_ac_read_mtp (
	.clk(clk),
	.d(\Selector23~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_mtp .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_mtp .power_up = "low";

cycloneiii_lcell_comb \sig_addr_cmd_state~40 (
	.dataa(\sig_addr_cmd_state~38_combout ),
	.datab(\sig_ac_req.s_ac_read_mtp~q ),
	.datac(\WideOr26~2_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~40_combout ),
	.cout());
defparam \sig_addr_cmd_state~40 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd_state~40 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_mtp (
	.clk(clk),
	.d(\sig_addr_cmd_state~40_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_mtp .power_up = "low";

cycloneiii_lcell_comb \ac_block:sig_count[7]~5 (
	.dataa(\ac_block:sig_count[7]~3_combout ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(\Equal13~1_combout ),
	.datad(\ac_block:sig_count[7]~4_combout ),
	.cin(gnd),
	.combout(\ac_block:sig_count[7]~5_combout ),
	.cout());
defparam \ac_block:sig_count[7]~5 .lut_mask = 16'hFEFF;
defparam \ac_block:sig_count[7]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector167~0 (
	.dataa(\ac_block:sig_count[7]~2_combout ),
	.datab(\Add23~12_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_count[7]~5_combout ),
	.cin(gnd),
	.combout(\Selector167~0_combout ),
	.cout());
defparam \Selector167~0 .lut_mask = 16'hEEFF;
defparam \Selector167~0 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[6] (
	.clk(clk),
	.d(\Selector167~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~7_combout ),
	.q(\ac_block:sig_count[6]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[6] .is_wysiwyg = "true";
defparam \ac_block:sig_count[6] .power_up = "low";

cycloneiii_lcell_comb \Selector170~1 (
	.dataa(\Selector170~0_combout ),
	.datab(\ac_block:sig_count[7]~2_combout ),
	.datac(\Add23~6_combout ),
	.datad(\ac_block:sig_count[7]~5_combout ),
	.cin(gnd),
	.combout(\Selector170~1_combout ),
	.cout());
defparam \Selector170~1 .lut_mask = 16'hFEFF;
defparam \Selector170~1 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[3] (
	.clk(clk),
	.d(\Selector170~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~7_combout ),
	.q(\ac_block:sig_count[3]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[3] .is_wysiwyg = "true";
defparam \ac_block:sig_count[3] .power_up = "low";

cycloneiii_lcell_comb \Selector171~0 (
	.dataa(\Add23~4_combout ),
	.datab(gnd),
	.datac(\ac_block:sig_count[1]~1_combout ),
	.datad(\ac_block:sig_count[7]~2_combout ),
	.cin(gnd),
	.combout(\Selector171~0_combout ),
	.cout());
defparam \Selector171~0 .lut_mask = 16'hAFFF;
defparam \Selector171~0 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[2] (
	.clk(clk),
	.d(\Selector171~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~7_combout ),
	.q(\ac_block:sig_count[2]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[2] .is_wysiwyg = "true";
defparam \ac_block:sig_count[2] .power_up = "low";

cycloneiii_lcell_comb \Selector175~3 (
	.dataa(\ac_block:sig_count[7]~q ),
	.datab(\ac_block:sig_count[6]~q ),
	.datac(\ac_block:sig_count[3]~q ),
	.datad(\ac_block:sig_count[2]~q ),
	.cin(gnd),
	.combout(\Selector175~3_combout ),
	.cout());
defparam \Selector175~3 .lut_mask = 16'h7FFF;
defparam \Selector175~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector175~4 (
	.dataa(\ac_block:sig_count[1]~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datad(\ac_block:sig_count[0]~q ),
	.cin(gnd),
	.combout(\Selector175~4_combout ),
	.cout());
defparam \Selector175~4 .lut_mask = 16'hFEFF;
defparam \Selector175~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector168~1 (
	.dataa(\ac_block:sig_count[7]~0_combout ),
	.datab(\Selector168~0_combout ),
	.datac(\Add23~10_combout ),
	.datad(\ac_block:sig_count[5]~2_combout ),
	.cin(gnd),
	.combout(\Selector168~1_combout ),
	.cout());
defparam \Selector168~1 .lut_mask = 16'hFAFC;
defparam \Selector168~1 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[5] (
	.clk(clk),
	.d(\Selector168~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[5]~4_combout ),
	.q(\ac_block:sig_count[5]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[5] .is_wysiwyg = "true";
defparam \ac_block:sig_count[5] .power_up = "low";

cycloneiii_lcell_comb \Selector169~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\Selector169~0_combout ),
	.cout());
defparam \Selector169~0 .lut_mask = 16'hEEFF;
defparam \Selector169~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_count~171 (
	.dataa(dgb_ac_access_gnt_r),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\sig_count~171_combout ),
	.cout());
defparam \sig_count~171 .lut_mask = 16'hAAFF;
defparam \sig_count~171 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector169~1_combout ),
	.cout());
defparam \Selector169~1 .lut_mask = 16'hEEEE;
defparam \Selector169~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~5 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(\Selector169~0_combout ),
	.datac(\sig_count~171_combout ),
	.datad(\Selector169~1_combout ),
	.cin(gnd),
	.combout(\Selector169~5_combout ),
	.cout());
defparam \Selector169~5 .lut_mask = 16'hFFFE;
defparam \Selector169~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~6 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datab(\Selector169~5_combout ),
	.datac(\ac_block:sig_burst_count[0]~q ),
	.datad(\Equal13~1_combout ),
	.cin(gnd),
	.combout(\Selector169~6_combout ),
	.cout());
defparam \Selector169~6 .lut_mask = 16'hEFFF;
defparam \Selector169~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector169~7 (
	.dataa(\Selector169~4_combout ),
	.datab(\Add23~8_combout ),
	.datac(\Selector169~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector169~7_combout ),
	.cout());
defparam \Selector169~7 .lut_mask = 16'hFEFE;
defparam \Selector169~7 .sum_lutc_input = "datac";

dffeas \ac_block:sig_count[4] (
	.clk(clk),
	.d(\Selector169~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_count[4]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[4] .is_wysiwyg = "true";
defparam \ac_block:sig_count[4] .power_up = "low";

cycloneiii_lcell_comb \Selector175~5 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\ac_block:sig_count[5]~q ),
	.datac(\ac_block:sig_count[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector175~5_combout ),
	.cout());
defparam \Selector175~5 .lut_mask = 16'hFEFE;
defparam \Selector175~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd_state~41 (
	.dataa(\sig_ac_req.s_ac_read_wd_lat~q ),
	.datab(\sig_addr_cmd_state~38_combout ),
	.datac(\WideOr26~2_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd_state~41_combout ),
	.cout());
defparam \sig_addr_cmd_state~41 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd_state~41 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat (
	.clk(clk),
	.d(\sig_addr_cmd_state~41_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat .power_up = "low";

cycloneiii_lcell_comb \Selector174~0 (
	.dataa(gnd),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.cin(gnd),
	.combout(\Selector174~0_combout ),
	.cout());
defparam \Selector174~0 .lut_mask = 16'h3FFF;
defparam \Selector174~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector174~1 (
	.dataa(\ac_block:sig_doing_rd_count~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(\Selector174~0_combout ),
	.datad(\dimm_driving_dq_proc~1_combout ),
	.cin(gnd),
	.combout(\Selector174~1_combout ),
	.cout());
defparam \Selector174~1 .lut_mask = 16'hEFFF;
defparam \Selector174~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector174~2 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector174~2_combout ),
	.cout());
defparam \Selector174~2 .lut_mask = 16'hEEEE;
defparam \Selector174~2 .sum_lutc_input = "datac";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat .power_up = "low";

cycloneiii_lcell_comb \Selector175~6 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(dgb_ac_access_gnt_r),
	.datac(\Equal13~1_combout ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.cin(gnd),
	.combout(\Selector175~6_combout ),
	.cout());
defparam \Selector175~6 .lut_mask = 16'hFFFE;
defparam \Selector175~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector175~7 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datac(\sig_dimm_driving_dq~q ),
	.datad(\Selector175~6_combout ),
	.cin(gnd),
	.combout(\Selector175~7_combout ),
	.cout());
defparam \Selector175~7 .lut_mask = 16'hFFEF;
defparam \Selector175~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector175~8 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\Selector174~1_combout ),
	.datac(\Selector174~2_combout ),
	.datad(\Selector175~7_combout ),
	.cin(gnd),
	.combout(\Selector175~8_combout ),
	.cout());
defparam \Selector175~8 .lut_mask = 16'hFFFD;
defparam \Selector175~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector175~9 (
	.dataa(\Selector175~3_combout ),
	.datab(\Selector175~4_combout ),
	.datac(\Selector175~5_combout ),
	.datad(\Selector175~8_combout ),
	.cin(gnd),
	.combout(\Selector175~9_combout ),
	.cout());
defparam \Selector175~9 .lut_mask = 16'hFFFE;
defparam \Selector175~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector165~0 (
	.dataa(\ac_block:sig_burst_count[0]~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datad(\Selector175~10_combout ),
	.cin(gnd),
	.combout(\Selector165~0_combout ),
	.cout());
defparam \Selector165~0 .lut_mask = 16'hBFFF;
defparam \Selector165~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal13~0 (
	.dataa(\Selector175~3_combout ),
	.datab(gnd),
	.datac(\ac_block:sig_count[5]~q ),
	.datad(\ac_block:sig_count[4]~q ),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'hAFFF;
defparam \Equal13~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector165~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datac(dgb_ac_access_gnt_r),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\Selector165~1_combout ),
	.cout());
defparam \Selector165~1 .lut_mask = 16'hFEFF;
defparam \Selector165~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector165~2 (
	.dataa(\Selector165~0_combout ),
	.datab(\Equal13~0_combout ),
	.datac(\Selector169~0_combout ),
	.datad(\Selector165~1_combout ),
	.cin(gnd),
	.combout(\Selector165~2_combout ),
	.cout());
defparam \Selector165~2 .lut_mask = 16'hFFFD;
defparam \Selector165~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector141~0 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(dgb_ac_access_gnt_r),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\Selector141~0_combout ),
	.cout());
defparam \Selector141~0 .lut_mask = 16'hEEFF;
defparam \Selector141~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector141~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.cin(gnd),
	.combout(\Selector141~1_combout ),
	.cout());
defparam \Selector141~1 .lut_mask = 16'hEEFF;
defparam \Selector141~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector141~2 (
	.dataa(\Selector138~0_combout ),
	.datab(\Selector141~0_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datad(\Selector141~1_combout ),
	.cin(gnd),
	.combout(\Selector141~2_combout ),
	.cout());
defparam \Selector141~2 .lut_mask = 16'hEFFF;
defparam \Selector141~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \btp_addr_array~0 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\btp_addr_array~0_combout ),
	.cout());
defparam \btp_addr_array~0 .lut_mask = 16'hEEEE;
defparam \btp_addr_array~0 .sum_lutc_input = "datac";

dffeas \ac_block:btp_addr_array[0][4] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btp_addr_array~0_combout ),
	.q(\ac_block:btp_addr_array[0][4]~q ),
	.prn(vcc));
defparam \ac_block:btp_addr_array[0][4] .is_wysiwyg = "true";
defparam \ac_block:btp_addr_array[0][4] .power_up = "low";

cycloneiii_lcell_comb \Selector141~3 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(\ac_block:btp_addr_array[0][4]~q ),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\Selector141~3_combout ),
	.cout());
defparam \Selector141~3 .lut_mask = 16'hFEFF;
defparam \Selector141~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector141~4 (
	.dataa(\Selector165~1_combout ),
	.datab(\ac_block:sig_count[0]~q ),
	.datac(\ac_block:sig_count[1]~q ),
	.datad(\Selector141~3_combout ),
	.cin(gnd),
	.combout(\Selector141~4_combout ),
	.cout());
defparam \Selector141~4 .lut_mask = 16'hFFBF;
defparam \Selector141~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector141~5 (
	.dataa(\Equal13~0_combout ),
	.datab(sig_addr_cmd0addr2),
	.datac(\Selector141~2_combout ),
	.datad(\Selector141~4_combout ),
	.cin(gnd),
	.combout(\Selector141~5_combout ),
	.cout());
defparam \Selector141~5 .lut_mask = 16'hFFEF;
defparam \Selector141~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd~435 (
	.dataa(\ac_block:sig_count[1]~q ),
	.datab(\Equal13~0_combout ),
	.datac(\ac_block:btp_addr_array[0][4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_addr_cmd~435_combout ),
	.cout());
defparam \sig_addr_cmd~435 .lut_mask = 16'hFEFE;
defparam \sig_addr_cmd~435 .sum_lutc_input = "datac";

dffeas \ctrl_dgrb_r.command_op.mtp_almt (
	.clk(clk),
	.d(\ctrl_dgrb.command_op.mtp_almt ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command_op.mtp_almt~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command_op.mtp_almt .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command_op.mtp_almt .power_up = "low";

dffeas current_mtp_almt(
	.clk(clk),
	.d(\ctrl_dgrb_r.command_op.mtp_almt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ac_muxctrl_broadcast_rcommand_req),
	.q(\current_mtp_almt~q ),
	.prn(vcc));
defparam current_mtp_almt.is_wysiwyg = "true";
defparam current_mtp_almt.power_up = "low";

dffeas \ac_block:btp_addr_array[0][3] (
	.clk(clk),
	.d(\current_mtp_almt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btp_addr_array~0_combout ),
	.q(\ac_block:btp_addr_array[0][3]~q ),
	.prn(vcc));
defparam \ac_block:btp_addr_array[0][3] .is_wysiwyg = "true";
defparam \ac_block:btp_addr_array[0][3] .power_up = "low";

cycloneiii_lcell_comb \Selector140~4 (
	.dataa(\Equal13~0_combout ),
	.datab(\ac_block:btp_addr_array[0][3]~q ),
	.datac(gnd),
	.datad(\ac_block:sig_count[1]~q ),
	.cin(gnd),
	.combout(\Selector140~4_combout ),
	.cout());
defparam \Selector140~4 .lut_mask = 16'hEEFF;
defparam \Selector140~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector140~5 (
	.dataa(\Selector169~0_combout ),
	.datab(\sig_addr_cmd~435_combout ),
	.datac(\Selector140~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector140~5_combout ),
	.cout());
defparam \Selector140~5 .lut_mask = 16'hFEFE;
defparam \Selector140~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector140~7 (
	.dataa(\Selector140~6_combout ),
	.datab(\Selector165~1_combout ),
	.datac(\Equal13~1_combout ),
	.datad(\current_mtp_almt~q ),
	.cin(gnd),
	.combout(\Selector140~7_combout ),
	.cout());
defparam \Selector140~7 .lut_mask = 16'hACFF;
defparam \Selector140~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector140~8 (
	.dataa(\Selector140~5_combout ),
	.datab(\Selector140~7_combout ),
	.datac(sig_addr_cmd0addr3),
	.datad(\Selector141~2_combout ),
	.cin(gnd),
	.combout(\Selector140~8_combout ),
	.cout());
defparam \Selector140~8 .lut_mask = 16'hFEFF;
defparam \Selector140~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~5 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(\Equal13~1_combout ),
	.datac(sig_addr_cmd0addr4),
	.datad(\Selector141~0_combout ),
	.cin(gnd),
	.combout(\Selector139~5_combout ),
	.cout());
defparam \Selector139~5 .lut_mask = 16'hFAFC;
defparam \Selector139~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd~436 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd~436_combout ),
	.cout());
defparam \sig_addr_cmd~436 .lut_mask = 16'hAAFF;
defparam \sig_addr_cmd~436 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~4 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.cin(gnd),
	.combout(\Selector139~4_combout ),
	.cout());
defparam \Selector139~4 .lut_mask = 16'hBFFF;
defparam \Selector139~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~9 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(\Selector139~4_combout ),
	.cin(gnd),
	.combout(\Selector139~9_combout ),
	.cout());
defparam \Selector139~9 .lut_mask = 16'hFDFF;
defparam \Selector139~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~6 (
	.dataa(sig_addr_cmd0addr4),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(\sig_addr_cmd~436_combout ),
	.datad(\Selector139~9_combout ),
	.cin(gnd),
	.combout(\Selector139~6_combout ),
	.cout());
defparam \Selector139~6 .lut_mask = 16'hFFFE;
defparam \Selector139~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~10 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(\ac_block:sig_burst_count[0]~q ),
	.datac(\ac_block:sig_count[1]~q ),
	.datad(\ac_block:btp_addr_array[0][4]~q ),
	.cin(gnd),
	.combout(\Selector139~10_combout ),
	.cout());
defparam \Selector139~10 .lut_mask = 16'hFFBF;
defparam \Selector139~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~7 (
	.dataa(\Equal13~0_combout ),
	.datab(sig_addr_cmd0addr4),
	.datac(\Selector139~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector139~7_combout ),
	.cout());
defparam \Selector139~7 .lut_mask = 16'hD8D8;
defparam \Selector139~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector139~8 (
	.dataa(\Selector139~5_combout ),
	.datab(\Selector139~6_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(\Selector139~7_combout ),
	.cin(gnd),
	.combout(\Selector139~8_combout ),
	.cout());
defparam \Selector139~8 .lut_mask = 16'hFFFE;
defparam \Selector139~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector138~1 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\Selector169~0_combout ),
	.datac(\sig_addr_cmd~435_combout ),
	.datad(\sig_addr_cmd~436_combout ),
	.cin(gnd),
	.combout(\Selector138~1_combout ),
	.cout());
defparam \Selector138~1 .lut_mask = 16'hFFFE;
defparam \Selector138~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector138~2 (
	.dataa(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datad(\sig_count~171_combout ),
	.cin(gnd),
	.combout(\Selector138~2_combout ),
	.cout());
defparam \Selector138~2 .lut_mask = 16'hEFFF;
defparam \Selector138~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd~434 (
	.dataa(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ac_block:sig_burst_count[0]~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd~434_combout ),
	.cout());
defparam \sig_addr_cmd~434 .lut_mask = 16'hAAFF;
defparam \sig_addr_cmd~434 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector140~9 (
	.dataa(\Selector175~3_combout ),
	.datab(\ac_block:sig_count[5]~q ),
	.datac(\ac_block:sig_count[4]~q ),
	.datad(\sig_addr_cmd~434_combout ),
	.cin(gnd),
	.combout(\Selector140~9_combout ),
	.cout());
defparam \Selector140~9 .lut_mask = 16'hFFBF;
defparam \Selector140~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector138~0 (
	.dataa(\Selector139~4_combout ),
	.datab(\Selector140~9_combout ),
	.datac(gnd),
	.datad(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.cin(gnd),
	.combout(\Selector138~0_combout ),
	.cout());
defparam \Selector138~0 .lut_mask = 16'hEEFF;
defparam \Selector138~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector138~3 (
	.dataa(\Selector138~1_combout ),
	.datab(sig_addr_cmd0addr5),
	.datac(\Selector138~2_combout ),
	.datad(\Selector138~0_combout ),
	.cin(gnd),
	.combout(\Selector138~3_combout ),
	.cout());
defparam \Selector138~3 .lut_mask = 16'hFEFF;
defparam \Selector138~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[12]~2 (
	.dataa(\sig_addr_cmd[0].addr[12]~1_combout ),
	.datab(\ac_block:sig_count[7]~0_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datad(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~2_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[12]~2 .lut_mask = 16'hACFF;
defparam \sig_addr_cmd[0].addr[12]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[12]~3 (
	.dataa(\sig_addr_cmd[0].addr[12]~0_combout ),
	.datab(\sig_addr_cmd[0].addr[12]~2_combout ),
	.datac(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(\Selector140~9_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~3_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[12]~3 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd[0].addr[12]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].cas_n~0 (
	.dataa(sig_addr_cmd0cas_n),
	.datab(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datac(gnd),
	.datad(\sig_addr_cmd[0].addr[12]~3_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].cas_n~0_combout ),
	.cout());
defparam \sig_addr_cmd[0].cas_n~0 .lut_mask = 16'hAACC;
defparam \sig_addr_cmd[0].cas_n~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_wd_lat~10 (
	.dataa(q_b_0),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_wd_lat~10_combout ),
	.cout());
defparam \sig_wd_lat~10 .lut_mask = 16'hEEEE;
defparam \sig_wd_lat~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgrb_main_block:sig_wd_lat[4]~0 (
	.dataa(\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(rdata_valid[0]),
	.datac(\sig_dimm_driving_dq~q ),
	.datad(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.cin(gnd),
	.combout(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.cout());
defparam \dgrb_main_block:sig_wd_lat[4]~0 .lut_mask = 16'hEFFF;
defparam \dgrb_main_block:sig_wd_lat[4]~0 .sum_lutc_input = "datac";

dffeas \dgrb_main_block:sig_wd_lat[0] (
	.clk(clk),
	.d(\sig_wd_lat~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[0]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[0] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[0] .power_up = "low";

cycloneiii_lcell_comb \wd_lat[0]~0 (
	.dataa(\dgrb_main_block:sig_wd_lat[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_lat[0]~0_combout ),
	.cout());
defparam \wd_lat[0]~0 .lut_mask = 16'h5555;
defparam \wd_lat[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_wd_lat~11 (
	.dataa(q_b_1),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_wd_lat~11_combout ),
	.cout());
defparam \sig_wd_lat~11 .lut_mask = 16'hEEEE;
defparam \sig_wd_lat~11 .sum_lutc_input = "datac";

dffeas \dgrb_main_block:sig_wd_lat[1] (
	.clk(clk),
	.d(\sig_wd_lat~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[1]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[1] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[1] .power_up = "low";

cycloneiii_lcell_comb \sig_wd_lat~12 (
	.dataa(q_b_4),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_wd_lat~12_combout ),
	.cout());
defparam \sig_wd_lat~12 .lut_mask = 16'hEEEE;
defparam \sig_wd_lat~12 .sum_lutc_input = "datac";

dffeas \dgrb_main_block:sig_wd_lat[4] (
	.clk(clk),
	.d(\sig_wd_lat~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[4]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[4] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[4] .power_up = "low";

cycloneiii_lcell_comb \sig_wd_lat~13 (
	.dataa(q_b_3),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_wd_lat~13_combout ),
	.cout());
defparam \sig_wd_lat~13 .lut_mask = 16'hEEEE;
defparam \sig_wd_lat~13 .sum_lutc_input = "datac";

dffeas \dgrb_main_block:sig_wd_lat[3] (
	.clk(clk),
	.d(\sig_wd_lat~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[3]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[3] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[3] .power_up = "low";

cycloneiii_lcell_comb \sig_wd_lat~14 (
	.dataa(q_b_2),
	.datab(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_wd_lat~14_combout ),
	.cout());
defparam \sig_wd_lat~14 .lut_mask = 16'hEEEE;
defparam \sig_wd_lat~14 .sum_lutc_input = "datac";

dffeas \dgrb_main_block:sig_wd_lat[2] (
	.clk(clk),
	.d(\sig_wd_lat~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[4]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[2]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[2] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[2] .power_up = "low";

cycloneiii_lcell_comb \wd_lat[2]~1 (
	.dataa(\dgrb_main_block:sig_wd_lat[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wd_lat[2]~1_combout ),
	.cout());
defparam \wd_lat[2]~1 .lut_mask = 16'h5555;
defparam \wd_lat[2]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_rdata_valid_lat_dec~3 (
	.dataa(rdata_valid[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dimm_driving_dq~q ),
	.cin(gnd),
	.combout(\seq_rdata_valid_lat_dec~3_combout ),
	.cout());
defparam \seq_rdata_valid_lat_dec~3 .lut_mask = 16'hAAFF;
defparam \seq_rdata_valid_lat_dec~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_rdata_valid_lat_dec~4 (
	.dataa(\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(\seq_rdata_valid_lat_dec~3_combout ),
	.datac(q_b_0),
	.datad(q_b_8),
	.cin(gnd),
	.combout(\seq_rdata_valid_lat_dec~4_combout ),
	.cout());
defparam \seq_rdata_valid_lat_dec~4 .lut_mask = 16'hFFFE;
defparam \seq_rdata_valid_lat_dec~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \pll_reconf_mux~1 (
	.dataa(\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(\sig_dgrb_state.s_reset_cdvw~q ),
	.datac(\sig_dgrb_state.s_test_phases~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pll_reconf_mux~1_combout ),
	.cout());
defparam \pll_reconf_mux~1 .lut_mask = 16'hFEFE;
defparam \pll_reconf_mux~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_pll_inc_dec_n~4 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_trk_pll_inc_dec_n~4_combout ),
	.cout());
defparam \sig_trk_pll_inc_dec_n~4 .lut_mask = 16'hEEEE;
defparam \sig_trk_pll_inc_dec_n~4 .sum_lutc_input = "datac";

dffeas \trk_block:sig_trk_last_state.s_trk_adjust_resync (
	.clk(clk),
	.d(\sig_trk_pll_inc_dec_n~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_adjust_resync .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_adjust_resync .power_up = "low";

cycloneiii_lcell_comb \sig_trk_pll_inc_dec_n~5 (
	.dataa(\LessThan10~2_combout ),
	.datab(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(\sig_trk_pll_inc_dec_n~q ),
	.datad(\sig_trk_pll_inc_dec_n~4_combout ),
	.cin(gnd),
	.combout(\sig_trk_pll_inc_dec_n~5_combout ),
	.cout());
defparam \sig_trk_pll_inc_dec_n~5 .lut_mask = 16'hF7D5;
defparam \sig_trk_pll_inc_dec_n~5 .sum_lutc_input = "datac";

dffeas sig_trk_pll_inc_dec_n(
	.clk(clk),
	.d(\sig_trk_pll_inc_dec_n~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_pll_inc_dec_n~q ),
	.prn(vcc));
defparam sig_trk_pll_inc_dec_n.is_wysiwyg = "true";
defparam sig_trk_pll_inc_dec_n.power_up = "low";

cycloneiii_lcell_comb \Add5~13 (
	.dataa(\Add5~6_combout ),
	.datab(\Add5~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~12 ),
	.combout(\Add5~13_combout ),
	.cout(\Add5~14 ));
defparam \Add5~13 .lut_mask = 16'h96BF;
defparam \Add5~13 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add5~15 (
	.dataa(\Add5~5_combout ),
	.datab(\Add5~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~14 ),
	.combout(\Add5~15_combout ),
	.cout(\Add5~16 ));
defparam \Add5~15 .lut_mask = 16'h96DF;
defparam \Add5~15 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add5~22 (
	.dataa(\Add9~8_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~17_combout ),
	.cin(gnd),
	.combout(\Add5~22_combout ),
	.cout());
defparam \Add5~22 .lut_mask = 16'h47FF;
defparam \Add5~22 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_num_phase_shifts[4] (
	.clk(clk),
	.d(\Add5~22_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[4]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[4] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[4] .power_up = "low";

cycloneiii_lcell_comb \Add5~23 (
	.dataa(\Add9~6_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~15_combout ),
	.cin(gnd),
	.combout(\Add5~23_combout ),
	.cout());
defparam \Add5~23 .lut_mask = 16'h47FF;
defparam \Add5~23 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_num_phase_shifts[3] (
	.clk(clk),
	.d(\Add5~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[3]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[3] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[3] .power_up = "low";

cycloneiii_lcell_comb \Add5~24 (
	.dataa(\Add9~4_combout ),
	.datab(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datac(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(\Add5~13_combout ),
	.cin(gnd),
	.combout(\Add5~24_combout ),
	.cout());
defparam \Add5~24 .lut_mask = 16'h47FF;
defparam \Add5~24 .sum_lutc_input = "datac";

dffeas \rsc_block:sig_num_phase_shifts[2] (
	.clk(clk),
	.d(\Add5~24_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_num_phase_shifts[2]~4_combout ),
	.q(\rsc_block:sig_num_phase_shifts[2]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[2] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[2] .power_up = "low";

cycloneiii_lcell_comb \Equal6~0 (
	.dataa(\rsc_block:sig_num_phase_shifts[5]~q ),
	.datab(\rsc_block:sig_num_phase_shifts[4]~q ),
	.datac(\rsc_block:sig_num_phase_shifts[3]~q ),
	.datad(\rsc_block:sig_num_phase_shifts[2]~q ),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h7FFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector59~0 (
	.dataa(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(\Equal6~0_combout ),
	.datac(\rsc_block:sig_num_phase_shifts[1]~q ),
	.datad(\rsc_block:sig_num_phase_shifts[0]~q ),
	.cin(gnd),
	.combout(\Selector59~0_combout ),
	.cout());
defparam \Selector59~0 .lut_mask = 16'hEFFF;
defparam \Selector59~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_rsc_pll_inc_dec_n~2 (
	.dataa(\rsc_block:sig_rewind_direction~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector59~0_combout ),
	.cin(gnd),
	.combout(\sig_rsc_pll_inc_dec_n~2_combout ),
	.cout());
defparam \sig_rsc_pll_inc_dec_n~2 .lut_mask = 16'hFF55;
defparam \sig_rsc_pll_inc_dec_n~2 .sum_lutc_input = "datac";

dffeas sig_rsc_pll_inc_dec_n(
	.clk(clk),
	.d(\sig_rsc_pll_inc_dec_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_pll_inc_dec_n~q ),
	.prn(vcc));
defparam sig_rsc_pll_inc_dec_n.is_wysiwyg = "true";
defparam sig_rsc_pll_inc_dec_n.power_up = "low";

cycloneiii_lcell_comb \seq_pll_inc_dec_n~2 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\pll_reconf_mux~1_combout ),
	.datac(\sig_trk_pll_inc_dec_n~q ),
	.datad(\sig_rsc_pll_inc_dec_n~q ),
	.cin(gnd),
	.combout(\seq_pll_inc_dec_n~2_combout ),
	.cout());
defparam \seq_pll_inc_dec_n~2 .lut_mask = 16'h8BFF;
defparam \seq_pll_inc_dec_n~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector59~2 (
	.dataa(\Selector59~1_combout ),
	.datab(\Selector59~0_combout ),
	.datac(\sig_phs_shft_busy~q ),
	.datad(\sig_phs_shft_busy_1t~q ),
	.cin(gnd),
	.combout(\Selector59~2_combout ),
	.cout());
defparam \Selector59~2 .lut_mask = 16'hEFFF;
defparam \Selector59~2 .sum_lutc_input = "datac";

dffeas sig_rsc_pll_start_reconfig(
	.clk(clk),
	.d(\Selector59~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_pll_start_reconfig~q ),
	.prn(vcc));
defparam sig_rsc_pll_start_reconfig.is_wysiwyg = "true";
defparam sig_rsc_pll_start_reconfig.power_up = "low";

cycloneiii_lcell_comb \Add16~0 (
	.dataa(\trk_block:sig_req_rsc_shift[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add16~0_combout ),
	.cout(\Add16~1 ));
defparam \Add16~0 .lut_mask = 16'hAA55;
defparam \Add16~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add16~14 (
	.dataa(\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add16~13 ),
	.combout(\Add16~14_combout ),
	.cout());
defparam \Add16~14 .lut_mask = 16'h5A5A;
defparam \Add16~14 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \sig_req_rsc_shift~66 (
	.dataa(\sig_req_rsc_shift~59_combout ),
	.datab(\Add16~14_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~66_combout ),
	.cout());
defparam \sig_req_rsc_shift~66 .lut_mask = 16'hEEFF;
defparam \sig_req_rsc_shift~66 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add17~1 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(gnd),
	.datac(gnd),
	.datad(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\Add17~1_combout ),
	.cout());
defparam \Add17~1 .lut_mask = 16'hAAFF;
defparam \Add17~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[5]~2 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datac(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datad(\Add17~1_combout ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[5]~2 .lut_mask = 16'hACFF;
defparam \trk_block:sig_req_rsc_shift[5]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~60 (
	.dataa(\trk_block:sig_mimic_cdv_found~q ),
	.datab(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~60_combout ),
	.cout());
defparam \sig_req_rsc_shift~60 .lut_mask = 16'hFEFF;
defparam \sig_req_rsc_shift~60 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~67 (
	.dataa(\sig_req_rsc_shift~65_combout ),
	.datab(\sig_req_rsc_shift~66_combout ),
	.datac(\sig_req_rsc_shift~60_combout ),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~67_combout ),
	.cout());
defparam \sig_req_rsc_shift~67 .lut_mask = 16'hFF7F;
defparam \sig_req_rsc_shift~67 .sum_lutc_input = "datac";

dffeas \trk_block:sig_req_rsc_shift[7] (
	.clk(clk),
	.d(\sig_req_rsc_shift~67_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_req_rsc_shift[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[7] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[7] .power_up = "low";

cycloneiii_lcell_comb \Add18~0 (
	.dataa(\trk_block:sig_req_rsc_shift[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add18~0_combout ),
	.cout(\Add18~1 ));
defparam \Add18~0 .lut_mask = 16'hAA55;
defparam \Add18~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Add18~2 (
	.dataa(\trk_block:sig_req_rsc_shift[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~1 ),
	.combout(\Add18~2_combout ),
	.cout(\Add18~3 ));
defparam \Add18~2 .lut_mask = 16'h5A5F;
defparam \Add18~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Add18~4 (
	.dataa(\trk_block:sig_req_rsc_shift[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add18~3 ),
	.combout(\Add18~4_combout ),
	.cout(\Add18~5 ));
defparam \Add18~4 .lut_mask = 16'h5AAF;
defparam \Add18~4 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[3]~0 (
	.dataa(\Add16~6_combout ),
	.datab(\Add18~6_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[3]~0_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[3]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_req_rsc_shift[3]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[2]~0 (
	.dataa(\Add16~4_combout ),
	.datab(\Add18~4_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[2]~0_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[2]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_req_rsc_shift[2]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[1]~0 (
	.dataa(\Add16~2_combout ),
	.datab(\Add18~2_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[1]~0_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[1]~0 .lut_mask = 16'hAACC;
defparam \trk_block:sig_req_rsc_shift[1]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~54 (
	.dataa(gnd),
	.datab(\trk_block:sig_req_rsc_shift[7]~q ),
	.datac(\LessThan10~1_combout ),
	.datad(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~54_combout ),
	.cout());
defparam \sig_req_rsc_shift~54 .lut_mask = 16'h3FFF;
defparam \sig_req_rsc_shift~54 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~55 (
	.dataa(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datab(\Add18~0_combout ),
	.datac(\Add16~0_combout ),
	.datad(\trk_block:sig_req_rsc_shift[7]~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~55_combout ),
	.cout());
defparam \sig_req_rsc_shift~55 .lut_mask = 16'hFAFC;
defparam \sig_req_rsc_shift~55 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~56 (
	.dataa(\Add15~0_combout ),
	.datab(\sig_req_rsc_shift~54_combout ),
	.datac(\sig_req_rsc_shift~55_combout ),
	.datad(\sig_trk_state~107_combout ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~56_combout ),
	.cout());
defparam \sig_req_rsc_shift~56 .lut_mask = 16'hFFFE;
defparam \sig_req_rsc_shift~56 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[5]~1 (
	.dataa(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datab(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(\trk_block:sig_req_rsc_shift[7]~q ),
	.datad(\LessThan10~1_combout ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[5]~1 .lut_mask = 16'hFFFE;
defparam \trk_block:sig_req_rsc_shift[5]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[5]~3 (
	.dataa(\trk_block:sig_mimic_cdv_found~q ),
	.datab(\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datac(gnd),
	.datad(\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[5]~3 .lut_mask = 16'hFF77;
defparam \trk_block:sig_req_rsc_shift[5]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_req_rsc_shift~57 (
	.dataa(\sig_dgrb_state.s_track~q ),
	.datab(\sig_req_rsc_shift~56_combout ),
	.datac(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datad(\trk_block:sig_req_rsc_shift[0]~q ),
	.cin(gnd),
	.combout(\sig_req_rsc_shift~57_combout ),
	.cout());
defparam \sig_req_rsc_shift~57 .lut_mask = 16'hFFF7;
defparam \sig_req_rsc_shift~57 .sum_lutc_input = "datac";

dffeas \trk_block:sig_req_rsc_shift[0] (
	.clk(clk),
	.d(\sig_req_rsc_shift~57_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_req_rsc_shift[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[0] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[0] .power_up = "low";

cycloneiii_lcell_comb \Add15~2 (
	.dataa(\trk_block:sig_mimic_delta[1]~q ),
	.datab(\trk_block:sig_req_rsc_shift[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~1 ),
	.combout(\Add15~2_combout ),
	.cout(\Add15~3 ));
defparam \Add15~2 .lut_mask = 16'h967F;
defparam \Add15~2 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \trk_block:sig_req_rsc_shift[5]~4 (
	.dataa(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datab(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(\sig_req_rsc_shift~54_combout ),
	.datad(\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.cin(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.cout());
defparam \trk_block:sig_req_rsc_shift[5]~4 .lut_mask = 16'h27FF;
defparam \trk_block:sig_req_rsc_shift[5]~4 .sum_lutc_input = "datac";

dffeas \trk_block:sig_req_rsc_shift[1] (
	.clk(clk),
	.d(\trk_block:sig_req_rsc_shift[1]~0_combout ),
	.asdata(\Add15~2_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sload(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.ena(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.q(\trk_block:sig_req_rsc_shift[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[1] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[1] .power_up = "low";

cycloneiii_lcell_comb \Add15~4 (
	.dataa(\trk_block:sig_mimic_delta[2]~q ),
	.datab(\trk_block:sig_req_rsc_shift[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add15~3 ),
	.combout(\Add15~4_combout ),
	.cout(\Add15~5 ));
defparam \Add15~4 .lut_mask = 16'h96EF;
defparam \Add15~4 .sum_lutc_input = "cin";

dffeas \trk_block:sig_req_rsc_shift[2] (
	.clk(clk),
	.d(\trk_block:sig_req_rsc_shift[2]~0_combout ),
	.asdata(\Add15~4_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sload(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.ena(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.q(\trk_block:sig_req_rsc_shift[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[2] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[2] .power_up = "low";

dffeas \trk_block:sig_req_rsc_shift[3] (
	.clk(clk),
	.d(\trk_block:sig_req_rsc_shift[3]~0_combout ),
	.asdata(\Add15~6_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sload(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.ena(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.q(\trk_block:sig_req_rsc_shift[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[3] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[3] .power_up = "low";

cycloneiii_lcell_comb \LessThan10~1 (
	.dataa(\LessThan10~0_combout ),
	.datab(\trk_block:sig_req_rsc_shift[3]~q ),
	.datac(\trk_block:sig_req_rsc_shift[2]~q ),
	.datad(\trk_block:sig_req_rsc_shift[1]~q ),
	.cin(gnd),
	.combout(\LessThan10~1_combout ),
	.cout());
defparam \LessThan10~1 .lut_mask = 16'hBFFF;
defparam \LessThan10~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_trk_state~106 (
	.dataa(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(gnd),
	.datac(\trk_block:sig_req_rsc_shift[7]~q ),
	.datad(\LessThan10~1_combout ),
	.cin(gnd),
	.combout(\sig_trk_state~106_combout ),
	.cout());
defparam \sig_trk_state~106 .lut_mask = 16'hAFFF;
defparam \sig_trk_state~106 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_phs_shft_start~0 (
	.dataa(\sig_phs_shft_busy~q ),
	.datab(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_phs_shft_start~0_combout ),
	.cout());
defparam \sig_phs_shft_start~0 .lut_mask = 16'hEEEE;
defparam \sig_phs_shft_start~0 .sum_lutc_input = "datac";

dffeas sig_phs_shft_start(
	.clk(clk),
	.d(\sig_phs_shft_start~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_start~q ),
	.prn(vcc));
defparam sig_phs_shft_start.is_wysiwyg = "true";
defparam sig_phs_shft_start.power_up = "low";

cycloneiii_lcell_comb \Selector126~0 (
	.dataa(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datab(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(\sig_trk_state~106_combout ),
	.datad(\sig_phs_shft_start~q ),
	.cin(gnd),
	.combout(\Selector126~0_combout ),
	.cout());
defparam \Selector126~0 .lut_mask = 16'hFEFF;
defparam \Selector126~0 .sum_lutc_input = "datac";

dffeas sig_trk_pll_start_reconfig(
	.clk(clk),
	.d(\Selector126~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_pll_start_reconfig~q ),
	.prn(vcc));
defparam sig_trk_pll_start_reconfig.is_wysiwyg = "true";
defparam sig_trk_pll_start_reconfig.power_up = "low";

cycloneiii_lcell_comb \seq_pll_start_reconfig~2 (
	.dataa(\sig_rsc_pll_start_reconfig~q ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\sig_trk_pll_start_reconfig~q ),
	.datad(\pll_reconf_mux~1_combout ),
	.cin(gnd),
	.combout(\seq_pll_start_reconfig~2_combout ),
	.cout());
defparam \seq_pll_start_reconfig~2 .lut_mask = 16'hFAFC;
defparam \seq_pll_start_reconfig~2 .sum_lutc_input = "datac";

dffeas \sig_dgrb_last_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgrb_state.s_release_admin~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_release_admin .power_up = "low";

cycloneiii_lcell_comb \ac_handshake_proc~1 (
	.dataa(\sig_dgrb_last_state.s_release_admin~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_idle~q ),
	.cin(gnd),
	.combout(\ac_handshake_proc~1_combout ),
	.cout());
defparam \ac_handshake_proc~1 .lut_mask = 16'hAAFF;
defparam \ac_handshake_proc~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_select~6 (
	.dataa(seq_ac_add_1t_ac_lat_internal),
	.datab(\pll_reconf_mux~1_combout ),
	.datac(gnd),
	.datad(\sig_dgrb_state.s_track~q ),
	.cin(gnd),
	.combout(\seq_pll_select~6_combout ),
	.cout());
defparam \seq_pll_select~6 .lut_mask = 16'hEEFF;
defparam \seq_pll_select~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \seq_pll_select~7 (
	.dataa(\pll_reconf_mux~1_combout ),
	.datab(\sig_dgrb_state.s_track~q ),
	.datac(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_pll_select~7_combout ),
	.cout());
defparam \seq_pll_select~7 .lut_mask = 16'hFEFE;
defparam \seq_pll_select~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~457 (
	.dataa(\sig_cdvw_state.current_window_size[5]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~457_combout ),
	.cout());
defparam \v_cdvw_state~457 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~457 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[5] (
	.clk(clk),
	.d(\v_cdvw_state~457_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[5] .power_up = "low";

cycloneiii_lcell_comb \dgrb_ctrl~8 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~8_combout ),
	.cout());
defparam \dgrb_ctrl~8 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~458 (
	.dataa(\sig_cdvw_state.current_window_size[4]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~458_combout ),
	.cout());
defparam \v_cdvw_state~458 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~458 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[4] (
	.clk(clk),
	.d(\v_cdvw_state~458_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[4] .power_up = "low";

cycloneiii_lcell_comb \dgrb_ctrl~9 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~9_combout ),
	.cout());
defparam \dgrb_ctrl~9 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~459 (
	.dataa(\sig_cdvw_state.current_window_size[3]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~459_combout ),
	.cout());
defparam \v_cdvw_state~459 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~459 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[3] (
	.clk(clk),
	.d(\v_cdvw_state~459_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[3] .power_up = "low";

cycloneiii_lcell_comb \dgrb_ctrl~10 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~10_combout ),
	.cout());
defparam \dgrb_ctrl~10 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \v_cdvw_state~460 (
	.dataa(\sig_cdvw_state.current_window_size[2]~q ),
	.datab(\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(\Selector32~0_combout ),
	.datad(\cdvw_proc~1_combout ),
	.cin(gnd),
	.combout(\v_cdvw_state~460_combout ),
	.cout());
defparam \v_cdvw_state~460 .lut_mask = 16'hEFFF;
defparam \v_cdvw_state~460 .sum_lutc_input = "datac";

dffeas \sig_cdvw_state.largest_window_size[2] (
	.clk(clk),
	.d(\v_cdvw_state~460_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.largest_window_size[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[2] .power_up = "low";

cycloneiii_lcell_comb \dgrb_ctrl~11 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~11_combout ),
	.cout());
defparam \dgrb_ctrl~11 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgrb_ctrl~12 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~12_combout ),
	.cout());
defparam \dgrb_ctrl~12 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgrb_ctrl~13 (
	.dataa(last_states_read_mtp),
	.datab(\sig_cdvw_state.largest_window_size[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgrb_ctrl~13_combout ),
	.cout());
defparam \dgrb_ctrl~13 .lut_mask = 16'hEEEE;
defparam \dgrb_ctrl~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_mmc_start~5 (
	.dataa(\trk_block:sig_trk_last_state.s_trk_mimic_sample~q ),
	.datab(\Equal10~0_combout ),
	.datac(\Equal10~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_mmc_start~5_combout ),
	.cout());
defparam \sig_mmc_start~5 .lut_mask = 16'h7F7F;
defparam \sig_mmc_start~5 .sum_lutc_input = "datac";

dffeas \trk_block:sig_mmc_start (
	.clk(clk),
	.d(\sig_mmc_start~5_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(vcc),
	.q(\trk_block:sig_mmc_start~q ),
	.prn(vcc));
defparam \trk_block:sig_mmc_start .is_wysiwyg = "true";
defparam \trk_block:sig_mmc_start .power_up = "low";

dffeas \trk_block:mimic_sample_req:v_echo (
	.clk(clk),
	.d(\trk_block:sig_mmc_start~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mimic_sample_req:v_echo~q ),
	.prn(vcc));
defparam \trk_block:mimic_sample_req:v_echo .is_wysiwyg = "true";
defparam \trk_block:mimic_sample_req:v_echo .power_up = "low";

cycloneiii_lcell_comb \seq_mmc_start~1 (
	.dataa(\trk_block:mimic_sample_req:v_echo~q ),
	.datab(\trk_block:sig_mmc_start~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\seq_mmc_start~1_combout ),
	.cout());
defparam \seq_mmc_start~1 .lut_mask = 16'hEEEE;
defparam \seq_mmc_start~1 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_dgwb (
	clk,
	sig_addr_cmd0addr2,
	sig_addr_cmd0addr3,
	sig_addr_cmd0addr4,
	sig_addr_cmd0addr5,
	sig_addr_cmd0cas_n,
	dgwb_wdata_24,
	dgwb_wdata_8,
	rst_n,
	dgwb_wdp_ovride1,
	dgwb_ac_access_req1,
	sig_addr_cmd0cs_n0,
	dgb_ac_access_gnt_r,
	ac_muxctrl_broadcast_rcommand_req,
	dgwb_ctrlcommand_done,
	curr_cmdcmd_write_btp,
	curr_cmdcmd_write_mtp,
	curr_cmdcmd_was,
	WideOr0,
	dgwb_wdata_25,
	dgwb_wdata_9,
	dgwb_wdata_26,
	dgwb_wdata_10,
	dgwb_wdata_27,
	dgwb_wdata_11,
	dgwb_wdata_28,
	dgwb_wdata_12,
	dgwb_wdata_29,
	dgwb_wdata_13,
	dgwb_wdata_30,
	dgwb_wdata_14,
	dgwb_wdata_31,
	dgwb_wdata_15)/* synthesis synthesis_greybox=1 */;
input 	clk;
output 	sig_addr_cmd0addr2;
output 	sig_addr_cmd0addr3;
output 	sig_addr_cmd0addr4;
output 	sig_addr_cmd0addr5;
output 	sig_addr_cmd0cas_n;
output 	dgwb_wdata_24;
output 	dgwb_wdata_8;
input 	rst_n;
output 	dgwb_wdp_ovride1;
output 	dgwb_ac_access_req1;
output 	sig_addr_cmd0cs_n0;
input 	dgb_ac_access_gnt_r;
input 	ac_muxctrl_broadcast_rcommand_req;
output 	dgwb_ctrlcommand_done;
input 	curr_cmdcmd_write_btp;
input 	curr_cmdcmd_write_mtp;
input 	curr_cmdcmd_was;
input 	WideOr0;
output 	dgwb_wdata_25;
output 	dgwb_wdata_9;
output 	dgwb_wdata_26;
output 	dgwb_wdata_10;
output 	dgwb_wdata_27;
output 	dgwb_wdata_11;
output 	dgwb_wdata_28;
output 	dgwb_wdata_12;
output 	dgwb_wdata_29;
output 	dgwb_wdata_13;
output 	dgwb_wdata_30;
output 	dgwb_wdata_14;
output 	dgwb_wdata_31;
output 	dgwb_wdata_15;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \Selector75~5_combout ;
wire \sig_dgwb_last_state.s_write_1100_step~q ;
wire \Selector50~1_combout ;
wire \Selector4~0_combout ;
wire \access_complete~q ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \Selector6~3_combout ;
wire \Selector7~0_combout ;
wire \Selector5~4_combout ;
wire \Selector5~5_combout ;
wire \Selector6~9_combout ;
wire \Selector12~2_combout ;
wire \Selector54~2_combout ;
wire \Selector75~7_combout ;
wire \Selector75~8_combout ;
wire \Selector75~9_combout ;
wire \Selector75~10_combout ;
wire \Selector13~0_combout ;
wire \sig_dgwb_state.s_release_admin~q ;
wire \sig_dgwb_state.s_idle~1_combout ;
wire \sig_dgwb_state.s_idle~q ;
wire \Selector4~1_combout ;
wire \sig_dgwb_state.s_wait_admin~q ;
wire \Selector6~4_combout ;
wire \Selector6~5_combout ;
wire \Selector5~2_combout ;
wire \sig_dgwb_state.s_write_btp~q ;
wire \Selector8~0_combout ;
wire \sig_dgwb_state.s_write_mtp~q ;
wire \Selector12~0_combout ;
wire \Selector6~6_combout ;
wire \Selector6~7_combout ;
wire \Selector11~0_combout ;
wire \sig_dgwb_state.s_write_0011_step~q ;
wire \ac_write_block:sig_count[0]~2 ;
wire \ac_write_block:sig_count[1]~2 ;
wire \ac_write_block:sig_count[2]~1_combout ;
wire \Selector6~8_combout ;
wire \sig_dgwb_state.s_write_ones~q ;
wire \sig_dgwb_last_state.s_write_ones~q ;
wire \Selector67~0_combout ;
wire \sig_dgwb_last_state.s_write_0011_step~q ;
wire \Selector10~1_combout ;
wire \sig_dgwb_state.s_write_1100_step~q ;
wire \Selector67~1_combout ;
wire \Selector7~1_combout ;
wire \Selector5~0_combout ;
wire \Selector12~1_combout ;
wire \Selector7~7_combout ;
wire \sig_dgwb_state.s_write_zeros~q ;
wire \Selector5~1_combout ;
wire \Selector5~8_combout ;
wire \sig_dgwb_last_state.s_write_01_pairs~q ;
wire \Selector10~0_combout ;
wire \Selector5~3_combout ;
wire \Selector5~9_combout ;
wire \Selector12~3_combout ;
wire \Selector12~4_combout ;
wire \sig_dgwb_state.s_write_wlat~q ;
wire \Selector7~2_combout ;
wire \sig_dgwb_last_state.s_write_wlat~q ;
wire \Selector5~6_combout ;
wire \Selector5~7_combout ;
wire \Selector7~3_combout ;
wire \Selector7~4_combout ;
wire \Selector7~5_combout ;
wire \Selector7~6_combout ;
wire \Selector9~0_combout ;
wire \sig_dgwb_state.s_write_01_pairs~q ;
wire \Selector67~2_combout ;
wire \Selector67~3_combout ;
wire \Selector67~4_combout ;
wire \sig_addr_cmd[0].addr[5]~1_combout ;
wire \generate_wdata~q ;
wire \ac_handshake_proc~11_combout ;
wire \ac_write_block:sig_count[2]~3_combout ;
wire \ac_write_block:sig_count[2]~q ;
wire \ac_write_block:sig_count[0]~1_combout ;
wire \ac_write_block:sig_count[0]~q ;
wire \ac_write_block:sig_count[1]~1_combout ;
wire \ac_write_block:sig_count[1]~q ;
wire \Selector75~6_combout ;
wire \ac_write_block:sig_count[2]~2 ;
wire \ac_write_block:sig_count[3]~2 ;
wire \ac_write_block:sig_count[4]~1_combout ;
wire \ac_write_block:sig_count[4]~q ;
wire \ac_write_block:sig_count[4]~2 ;
wire \ac_write_block:sig_count[5]~2 ;
wire \ac_write_block:sig_count[6]~1_combout ;
wire \ac_write_block:sig_count[6]~q ;
wire \Equal1~0_combout ;
wire \Equal0~0_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \sig_addr_cmd[0].addr[5]~0_combout ;
wire \sig_dgwb_last_state.s_write_zeros~q ;
wire \sig_addr_cmd[0].addr[5]~2_combout ;
wire \sig_addr_cmd[0].addr[5]~3_combout ;
wire \sig_addr_cmd[0].addr[5]~4_combout ;
wire \sig_addr_cmd[0].addr[5]~5_combout ;
wire \sig_addr_cmd~518_combout ;
wire \Equal4~0_combout ;
wire \sig_addr_cmd[0].addr[5]~6_combout ;
wire \sig_addr_cmd[0].addr[5]~7_combout ;
wire \Selector25~0_combout ;
wire \ac_write_block:sig_count[3]~1_combout ;
wire \ac_write_block:sig_count[3]~q ;
wire \Equal1~1_combout ;
wire \Selector24~0_combout ;
wire \Selector23~0_combout ;
wire \Selector58~0_combout ;
wire \dgwb_wdata[24]~9_combout ;
wire \dgwb_wdata~11_combout ;
wire \Selector66~0_combout ;
wire \dgwb_wdata[8]~10_combout ;
wire \dgwb_dqs_burst~0_combout ;
wire \Selector6~0_combout ;
wire \Selector50~0_combout ;
wire \Selector50~2_combout ;
wire \Selector50~3_combout ;
wire \sig_dgwb_last_state.s_release_admin~q ;
wire \ac_handshake_proc~2_combout ;
wire \Selector57~0_combout ;
wire \Selector65~0_combout ;
wire \Selector56~0_combout ;
wire \Selector64~0_combout ;
wire \Selector55~0_combout ;
wire \Selector63~0_combout ;
wire \Selector54~3_combout ;
wire \Selector62~2_combout ;
wire \ac_write_block:sig_count[5]~1_combout ;
wire \ac_write_block:sig_count[5]~q ;
wire \Selector53~0_combout ;
wire \Selector61~0_combout ;
wire \Selector52~0_combout ;
wire \Selector60~0_combout ;
wire \ac_write_block:sig_count[6]~2 ;
wire \ac_write_block:sig_count[7]~1_combout ;
wire \ac_write_block:sig_count[7]~q ;
wire \Selector51~0_combout ;
wire \Selector59~0_combout ;


cycloneiii_lcell_comb \Selector75~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_write_block:sig_count[5]~q ),
	.datad(\ac_write_block:sig_count[7]~q ),
	.cin(gnd),
	.combout(\Selector75~5_combout ),
	.cout());
defparam \Selector75~5 .lut_mask = 16'h0FFF;
defparam \Selector75~5 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_write_1100_step (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_1100_step~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_1100_step~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_1100_step .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_1100_step .power_up = "low";

cycloneiii_lcell_comb \Selector50~1 (
	.dataa(\sig_dgwb_last_state.s_write_1100_step~q ),
	.datab(\sig_dgwb_last_state.s_write_0011_step~q ),
	.datac(\sig_dgwb_state.s_write_0011_step~q ),
	.datad(\sig_dgwb_state.s_write_1100_step~q ),
	.cin(gnd),
	.combout(\Selector50~1_combout ),
	.cout());
defparam \Selector50~1 .lut_mask = 16'hEFFF;
defparam \Selector50~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector4~0 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(WideOr0),
	.datac(gnd),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hEEFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas access_complete(
	.clk(clk),
	.d(\Selector75~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\access_complete~q ),
	.prn(vcc));
defparam access_complete.is_wysiwyg = "true";
defparam access_complete.power_up = "low";

cycloneiii_lcell_comb \Selector6~1 (
	.dataa(\sig_dgwb_last_state.s_write_wlat~q ),
	.datab(\sig_dgwb_last_state.s_write_0011_step~q ),
	.datac(\sig_dgwb_state.s_write_0011_step~q ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hFAFC;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~2 (
	.dataa(\access_complete~q ),
	.datab(\sig_dgwb_last_state.s_write_ones~q ),
	.datac(\Selector6~1_combout ),
	.datad(\sig_dgwb_state.s_write_ones~q ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hFAFC;
defparam \Selector6~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~3 (
	.dataa(\access_complete~q ),
	.datab(\Selector6~0_combout ),
	.datac(\Selector10~0_combout ),
	.datad(\sig_addr_cmd[0].addr[5]~4_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
defparam \Selector6~3 .lut_mask = 16'hFFFE;
defparam \Selector6~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~0 (
	.dataa(\sig_dgwb_state.s_write_btp~q ),
	.datab(\sig_dgwb_state.s_wait_admin~q ),
	.datac(gnd),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hEEFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~4 (
	.dataa(\sig_dgwb_state.s_write_ones~q ),
	.datab(\sig_dgwb_last_state.s_write_ones~q ),
	.datac(\access_complete~q ),
	.datad(\sig_dgwb_state.s_write_zeros~q ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
defparam \Selector5~4 .lut_mask = 16'hFEFF;
defparam \Selector5~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~5 (
	.dataa(\sig_dgwb_last_state.s_write_1100_step~q ),
	.datab(\sig_dgwb_last_state.s_write_0011_step~q ),
	.datac(\sig_dgwb_state.s_write_0011_step~q ),
	.datad(\sig_dgwb_state.s_write_1100_step~q ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
defparam \Selector5~5 .lut_mask = 16'hFAFC;
defparam \Selector5~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~9 (
	.dataa(\sig_dgwb_state.s_write_zeros~q ),
	.datab(\sig_dgwb_last_state.s_write_zeros~q ),
	.datac(\access_complete~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector6~9_combout ),
	.cout());
defparam \Selector6~9 .lut_mask = 16'hFEFE;
defparam \Selector6~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~2 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(\Selector12~0_combout ),
	.datac(dgb_ac_access_gnt_r),
	.datad(curr_cmdcmd_was),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
defparam \Selector12~2 .lut_mask = 16'hFFFE;
defparam \Selector12~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector54~2 (
	.dataa(\ac_write_block:sig_count[4]~q ),
	.datab(\sig_dgwb_state.s_write_wlat~q ),
	.datac(\generate_wdata~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector54~2_combout ),
	.cout());
defparam \Selector54~2 .lut_mask = 16'hFEFE;
defparam \Selector54~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector75~7 (
	.dataa(\Selector75~6_combout ),
	.datab(\Selector54~2_combout ),
	.datac(\ac_write_block:sig_count[3]~q ),
	.datad(\ac_write_block:sig_count[2]~q ),
	.cin(gnd),
	.combout(\Selector75~7_combout ),
	.cout());
defparam \Selector75~7 .lut_mask = 16'hEFFF;
defparam \Selector75~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector75~8 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\ac_write_block:sig_count[2]~q ),
	.datac(\ac_write_block:sig_count[0]~q ),
	.datad(\ac_write_block:sig_count[4]~q ),
	.cin(gnd),
	.combout(\Selector75~8_combout ),
	.cout());
defparam \Selector75~8 .lut_mask = 16'hFEFF;
defparam \Selector75~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector75~9 (
	.dataa(\ac_write_block:sig_count[1]~q ),
	.datab(\Selector75~8_combout ),
	.datac(gnd),
	.datad(\Selector5~1_combout ),
	.cin(gnd),
	.combout(\Selector75~9_combout ),
	.cout());
defparam \Selector75~9 .lut_mask = 16'hFFEE;
defparam \Selector75~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector75~10 (
	.dataa(\Selector75~5_combout ),
	.datab(\ac_write_block:sig_count[6]~q ),
	.datac(\Selector75~7_combout ),
	.datad(\Selector75~9_combout ),
	.cin(gnd),
	.combout(\Selector75~10_combout ),
	.cout());
defparam \Selector75~10 .lut_mask = 16'hFFFE;
defparam \Selector75~10 .sum_lutc_input = "datac";

dffeas \sig_addr_cmd[0].addr[2] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dgwb_state.s_write_wlat~q ),
	.sload(\sig_dgwb_state.s_write_1100_step~q ),
	.ena(\sig_addr_cmd[0].addr[5]~7_combout ),
	.q(sig_addr_cmd0addr2),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[2] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[2] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[3] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dgwb_state.s_write_wlat~q ),
	.sload(\sig_dgwb_state.s_write_1100_step~q ),
	.ena(\sig_addr_cmd[0].addr[5]~7_combout ),
	.q(sig_addr_cmd0addr3),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[3] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[3] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[4] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[5]~7_combout ),
	.q(sig_addr_cmd0addr4),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[4] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[4] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[5] (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[5]~7_combout ),
	.q(sig_addr_cmd0addr5),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[5] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[5] .power_up = "low";

dffeas \sig_addr_cmd[0].cas_n (
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[5]~7_combout ),
	.q(sig_addr_cmd0cas_n),
	.prn(vcc));
defparam \sig_addr_cmd[0].cas_n .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cas_n .power_up = "low";

dffeas \dgwb_wdata[24] (
	.clk(clk),
	.d(\dgwb_wdata[24]~9_combout ),
	.asdata(\dgwb_wdata~11_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(vcc),
	.q(dgwb_wdata_24),
	.prn(vcc));
defparam \dgwb_wdata[24] .is_wysiwyg = "true";
defparam \dgwb_wdata[24] .power_up = "low";

dffeas \dgwb_wdata[8] (
	.clk(clk),
	.d(\dgwb_wdata[8]~10_combout ),
	.asdata(\dgwb_wdata~11_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(vcc),
	.q(dgwb_wdata_8),
	.prn(vcc));
defparam \dgwb_wdata[8] .is_wysiwyg = "true";
defparam \dgwb_wdata[8] .power_up = "low";

dffeas dgwb_wdp_ovride(
	.clk(clk),
	.d(\dgwb_dqs_burst~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdp_ovride1),
	.prn(vcc));
defparam dgwb_wdp_ovride.is_wysiwyg = "true";
defparam dgwb_wdp_ovride.power_up = "low";

dffeas dgwb_ac_access_req(
	.clk(clk),
	.d(\ac_handshake_proc~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_ac_access_req1),
	.prn(vcc));
defparam dgwb_ac_access_req.is_wysiwyg = "true";
defparam dgwb_ac_access_req.power_up = "low";

dffeas \sig_addr_cmd[0].cs_n[0] (
	.clk(clk),
	.d(\Selector50~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0cs_n0),
	.prn(vcc));
defparam \sig_addr_cmd[0].cs_n[0] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cs_n[0] .power_up = "low";

dffeas \dgwb_ctrl.command_done (
	.clk(clk),
	.d(\ac_handshake_proc~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_ctrlcommand_done),
	.prn(vcc));
defparam \dgwb_ctrl.command_done .is_wysiwyg = "true";
defparam \dgwb_ctrl.command_done .power_up = "low";

dffeas \dgwb_wdata[25] (
	.clk(clk),
	.d(\Selector57~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_25),
	.prn(vcc));
defparam \dgwb_wdata[25] .is_wysiwyg = "true";
defparam \dgwb_wdata[25] .power_up = "low";

dffeas \dgwb_wdata[9] (
	.clk(clk),
	.d(\Selector65~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_9),
	.prn(vcc));
defparam \dgwb_wdata[9] .is_wysiwyg = "true";
defparam \dgwb_wdata[9] .power_up = "low";

dffeas \dgwb_wdata[26] (
	.clk(clk),
	.d(\Selector56~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_26),
	.prn(vcc));
defparam \dgwb_wdata[26] .is_wysiwyg = "true";
defparam \dgwb_wdata[26] .power_up = "low";

dffeas \dgwb_wdata[10] (
	.clk(clk),
	.d(\Selector64~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_10),
	.prn(vcc));
defparam \dgwb_wdata[10] .is_wysiwyg = "true";
defparam \dgwb_wdata[10] .power_up = "low";

dffeas \dgwb_wdata[27] (
	.clk(clk),
	.d(\Selector55~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_27),
	.prn(vcc));
defparam \dgwb_wdata[27] .is_wysiwyg = "true";
defparam \dgwb_wdata[27] .power_up = "low";

dffeas \dgwb_wdata[11] (
	.clk(clk),
	.d(\Selector63~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_11),
	.prn(vcc));
defparam \dgwb_wdata[11] .is_wysiwyg = "true";
defparam \dgwb_wdata[11] .power_up = "low";

dffeas \dgwb_wdata[28] (
	.clk(clk),
	.d(\Selector54~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_28),
	.prn(vcc));
defparam \dgwb_wdata[28] .is_wysiwyg = "true";
defparam \dgwb_wdata[28] .power_up = "low";

dffeas \dgwb_wdata[12] (
	.clk(clk),
	.d(\Selector62~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_12),
	.prn(vcc));
defparam \dgwb_wdata[12] .is_wysiwyg = "true";
defparam \dgwb_wdata[12] .power_up = "low";

dffeas \dgwb_wdata[29] (
	.clk(clk),
	.d(\Selector53~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_29),
	.prn(vcc));
defparam \dgwb_wdata[29] .is_wysiwyg = "true";
defparam \dgwb_wdata[29] .power_up = "low";

dffeas \dgwb_wdata[13] (
	.clk(clk),
	.d(\Selector61~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_13),
	.prn(vcc));
defparam \dgwb_wdata[13] .is_wysiwyg = "true";
defparam \dgwb_wdata[13] .power_up = "low";

dffeas \dgwb_wdata[30] (
	.clk(clk),
	.d(\Selector52~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_30),
	.prn(vcc));
defparam \dgwb_wdata[30] .is_wysiwyg = "true";
defparam \dgwb_wdata[30] .power_up = "low";

dffeas \dgwb_wdata[14] (
	.clk(clk),
	.d(\Selector60~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_14),
	.prn(vcc));
defparam \dgwb_wdata[14] .is_wysiwyg = "true";
defparam \dgwb_wdata[14] .power_up = "low";

dffeas \dgwb_wdata[31] (
	.clk(clk),
	.d(\Selector51~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_31),
	.prn(vcc));
defparam \dgwb_wdata[31] .is_wysiwyg = "true";
defparam \dgwb_wdata[31] .power_up = "low";

dffeas \dgwb_wdata[15] (
	.clk(clk),
	.d(\Selector59~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_15),
	.prn(vcc));
defparam \dgwb_wdata[15] .is_wysiwyg = "true";
defparam \dgwb_wdata[15] .power_up = "low";

cycloneiii_lcell_comb \Selector13~0 (
	.dataa(\Selector6~2_combout ),
	.datab(dgb_ac_access_gnt_r),
	.datac(\sig_dgwb_state.s_release_admin~q ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hEFFE;
defparam \Selector13~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_release_admin (
	.clk(clk),
	.d(\Selector13~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_release_admin .power_up = "low";

cycloneiii_lcell_comb \sig_dgwb_state.s_idle~1 (
	.dataa(dgb_ac_access_gnt_r),
	.datab(\sig_dgwb_state.s_idle~q ),
	.datac(\Selector6~6_combout ),
	.datad(\sig_dgwb_state.s_release_admin~q ),
	.cin(gnd),
	.combout(\sig_dgwb_state.s_idle~1_combout ),
	.cout());
defparam \sig_dgwb_state.s_idle~1 .lut_mask = 16'hACFF;
defparam \sig_dgwb_state.s_idle~1 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_idle (
	.clk(clk),
	.d(\sig_dgwb_state.s_idle~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_idle .power_up = "low";

cycloneiii_lcell_comb \Selector4~1 (
	.dataa(\Selector4~0_combout ),
	.datab(ac_muxctrl_broadcast_rcommand_req),
	.datac(\sig_dgwb_state.s_idle~q ),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hEFFF;
defparam \Selector4~1 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_wait_admin (
	.clk(clk),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_wait_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_wait_admin .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_wait_admin .power_up = "low";

cycloneiii_lcell_comb \Selector6~4 (
	.dataa(\Selector6~3_combout ),
	.datab(\sig_dgwb_state.s_wait_admin~q ),
	.datac(\sig_dgwb_state.s_release_admin~q ),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
defparam \Selector6~4 .lut_mask = 16'hFEFF;
defparam \Selector6~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~5 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(ac_muxctrl_broadcast_rcommand_req),
	.datac(\sig_dgwb_state.s_idle~q ),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
defparam \Selector6~5 .lut_mask = 16'hEFFF;
defparam \Selector6~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~2 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(dgb_ac_access_gnt_r),
	.datac(curr_cmdcmd_write_btp),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hFEFE;
defparam \Selector5~2 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_btp (
	.clk(clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_btp~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_btp .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_btp .power_up = "low";

cycloneiii_lcell_comb \Selector8~0 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(dgb_ac_access_gnt_r),
	.datac(curr_cmdcmd_write_mtp),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFEFE;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_mtp (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_mtp~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_mtp .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_mtp .power_up = "low";

cycloneiii_lcell_comb \Selector12~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sig_dgwb_state.s_write_btp~q ),
	.datad(\sig_dgwb_state.s_write_mtp~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'h0FFF;
defparam \Selector12~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~6 (
	.dataa(\Selector6~2_combout ),
	.datab(\Selector6~4_combout ),
	.datac(\Selector6~5_combout ),
	.datad(\Selector12~0_combout ),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
defparam \Selector6~6 .lut_mask = 16'hFEFF;
defparam \Selector6~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~7 (
	.dataa(\access_complete~q ),
	.datab(\Selector6~6_combout ),
	.datac(dgb_ac_access_gnt_r),
	.datad(\sig_dgwb_state.s_release_admin~q ),
	.cin(gnd),
	.combout(\Selector6~7_combout ),
	.cout());
defparam \Selector6~7 .lut_mask = 16'hFEFF;
defparam \Selector6~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector11~0 (
	.dataa(\sig_addr_cmd[0].addr[5]~4_combout ),
	.datab(\Selector6~7_combout ),
	.datac(\sig_dgwb_state.s_write_0011_step~q ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'hFEFF;
defparam \Selector11~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_0011_step (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_0011_step~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_0011_step .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_0011_step .power_up = "low";

cycloneiii_lcell_comb \ac_write_block:sig_count[0]~1 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ac_write_block:sig_count[0]~1_combout ),
	.cout(\ac_write_block:sig_count[0]~2 ));
defparam \ac_write_block:sig_count[0]~1 .lut_mask = 16'h55AA;
defparam \ac_write_block:sig_count[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_write_block:sig_count[1]~1 (
	.dataa(\ac_write_block:sig_count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[0]~2 ),
	.combout(\ac_write_block:sig_count[1]~1_combout ),
	.cout(\ac_write_block:sig_count[1]~2 ));
defparam \ac_write_block:sig_count[1]~1 .lut_mask = 16'h5A5F;
defparam \ac_write_block:sig_count[1]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \ac_write_block:sig_count[2]~1 (
	.dataa(\ac_write_block:sig_count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[1]~2 ),
	.combout(\ac_write_block:sig_count[2]~1_combout ),
	.cout(\ac_write_block:sig_count[2]~2 ));
defparam \ac_write_block:sig_count[2]~1 .lut_mask = 16'h5AAF;
defparam \ac_write_block:sig_count[2]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \Selector6~8 (
	.dataa(\Selector6~0_combout ),
	.datab(\Selector6~7_combout ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(\Selector6~8_combout ),
	.cout());
defparam \Selector6~8 .lut_mask = 16'hFEFF;
defparam \Selector6~8 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_ones (
	.clk(clk),
	.d(\Selector6~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_ones~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_ones .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_ones .power_up = "low";

dffeas \sig_dgwb_last_state.s_write_ones (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_ones~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_ones~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_ones .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_ones .power_up = "low";

cycloneiii_lcell_comb \Selector67~0 (
	.dataa(\sig_dgwb_state.s_write_ones~q ),
	.datab(\sig_dgwb_last_state.s_write_ones~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector67~0_combout ),
	.cout());
defparam \Selector67~0 .lut_mask = 16'hEEEE;
defparam \Selector67~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_write_0011_step (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_0011_step~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_0011_step~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_0011_step .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_0011_step .power_up = "low";

cycloneiii_lcell_comb \Selector10~1 (
	.dataa(\Selector10~0_combout ),
	.datab(\Selector6~7_combout ),
	.datac(\sig_dgwb_state.s_write_1100_step~q ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hFEFF;
defparam \Selector10~1 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_1100_step (
	.clk(clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_1100_step~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_1100_step .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_1100_step .power_up = "low";

cycloneiii_lcell_comb \Selector67~1 (
	.dataa(\sig_dgwb_last_state.s_write_1100_step~q ),
	.datab(\sig_dgwb_last_state.s_write_0011_step~q ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_1100_step~q ),
	.cin(gnd),
	.combout(\Selector67~1_combout ),
	.cout());
defparam \Selector67~1 .lut_mask = 16'hAACC;
defparam \Selector67~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~1 (
	.dataa(\sig_dgwb_state.s_idle~q ),
	.datab(ac_muxctrl_broadcast_rcommand_req),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_mtp~q ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'hEEFF;
defparam \Selector7~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sig_dgwb_state.s_write_1100_step~q ),
	.datad(\sig_dgwb_state.s_write_0011_step~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'h0FFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~1 (
	.dataa(gnd),
	.datab(\sig_dgwb_state.s_wait_admin~q ),
	.datac(\sig_dgwb_state.s_write_btp~q ),
	.datad(\sig_dgwb_state.s_write_mtp~q ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
defparam \Selector12~1 .lut_mask = 16'h3FFF;
defparam \Selector12~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~7 (
	.dataa(\sig_dgwb_state.s_write_btp~q ),
	.datab(\sig_dgwb_state.s_write_zeros~q ),
	.datac(\Selector7~6_combout ),
	.datad(\sig_dgwb_state.s_write_mtp~q ),
	.cin(gnd),
	.combout(\Selector7~7_combout ),
	.cout());
defparam \Selector7~7 .lut_mask = 16'hEFFF;
defparam \Selector7~7 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_zeros (
	.clk(clk),
	.d(\Selector7~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_zeros~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_zeros .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_zeros .power_up = "low";

cycloneiii_lcell_comb \Selector5~1 (
	.dataa(\Selector5~0_combout ),
	.datab(\sig_dgwb_state.s_write_zeros~q ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\sig_dgwb_state.s_write_01_pairs~q ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFFFD;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~8 (
	.dataa(\Selector6~9_combout ),
	.datab(\sig_dgwb_state.s_release_admin~q ),
	.datac(\Selector5~1_combout ),
	.datad(dgb_ac_access_gnt_r),
	.cin(gnd),
	.combout(\Selector5~8_combout ),
	.cout());
defparam \Selector5~8 .lut_mask = 16'hEFFF;
defparam \Selector5~8 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_write_01_pairs (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_01_pairs~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_01_pairs~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_01_pairs .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_01_pairs .power_up = "low";

cycloneiii_lcell_comb \Selector10~0 (
	.dataa(\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hEEEE;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~3 (
	.dataa(\access_complete~q ),
	.datab(gnd),
	.datac(\sig_dgwb_state.s_write_zeros~q ),
	.datad(\sig_dgwb_state.s_write_ones~q ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
defparam \Selector5~3 .lut_mask = 16'hAFFF;
defparam \Selector5~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~9 (
	.dataa(\Selector5~7_combout ),
	.datab(\Selector5~8_combout ),
	.datac(\Selector10~0_combout ),
	.datad(\Selector5~3_combout ),
	.cin(gnd),
	.combout(\Selector5~9_combout ),
	.cout());
defparam \Selector5~9 .lut_mask = 16'hFFFE;
defparam \Selector5~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~3 (
	.dataa(WideOr0),
	.datab(ac_muxctrl_broadcast_rcommand_req),
	.datac(\sig_dgwb_state.s_idle~q ),
	.datad(\Selector5~9_combout ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
defparam \Selector12~3 .lut_mask = 16'hA3FF;
defparam \Selector12~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector12~4 (
	.dataa(\Selector12~2_combout ),
	.datab(\Selector12~1_combout ),
	.datac(\sig_dgwb_state.s_write_wlat~q ),
	.datad(\Selector12~3_combout ),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
defparam \Selector12~4 .lut_mask = 16'hFFFE;
defparam \Selector12~4 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_wlat (
	.clk(clk),
	.d(\Selector12~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_wlat~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_wlat .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_wlat .power_up = "low";

cycloneiii_lcell_comb \Selector7~2 (
	.dataa(\sig_dgwb_state.s_write_ones~q ),
	.datab(\sig_dgwb_state.s_release_admin~q ),
	.datac(\sig_dgwb_state.s_write_wlat~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector7~2_combout ),
	.cout());
defparam \Selector7~2 .lut_mask = 16'hFEFE;
defparam \Selector7~2 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_write_wlat (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_wlat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_wlat~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_wlat .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_wlat .power_up = "low";

cycloneiii_lcell_comb \Selector5~6 (
	.dataa(\Selector5~5_combout ),
	.datab(\sig_dgwb_last_state.s_write_wlat~q ),
	.datac(\Selector5~0_combout ),
	.datad(\sig_dgwb_state.s_release_admin~q ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
defparam \Selector5~6 .lut_mask = 16'hFEFF;
defparam \Selector5~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector5~7 (
	.dataa(\Selector5~4_combout ),
	.datab(\Selector5~6_combout ),
	.datac(\Selector5~3_combout ),
	.datad(\sig_dgwb_state.s_write_01_pairs~q ),
	.cin(gnd),
	.combout(\Selector5~7_combout ),
	.cout());
defparam \Selector5~7 .lut_mask = 16'hFEFF;
defparam \Selector5~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~3 (
	.dataa(\Selector10~0_combout ),
	.datab(\Selector5~3_combout ),
	.datac(\Selector5~7_combout ),
	.datad(\Selector5~8_combout ),
	.cin(gnd),
	.combout(\Selector7~3_combout ),
	.cout());
defparam \Selector7~3 .lut_mask = 16'hFFFE;
defparam \Selector7~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~4 (
	.dataa(\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(\Selector5~0_combout ),
	.datac(\Selector7~2_combout ),
	.datad(\Selector7~3_combout ),
	.cin(gnd),
	.combout(\Selector7~4_combout ),
	.cout());
defparam \Selector7~4 .lut_mask = 16'hFFFB;
defparam \Selector7~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~5 (
	.dataa(\Selector6~9_combout ),
	.datab(\sig_dgwb_state.s_wait_admin~q ),
	.datac(\sig_dgwb_state.s_idle~q ),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector7~5_combout ),
	.cout());
defparam \Selector7~5 .lut_mask = 16'hEFFF;
defparam \Selector7~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector7~6 (
	.dataa(\Selector7~0_combout ),
	.datab(\Selector7~1_combout ),
	.datac(\Selector7~4_combout ),
	.datad(\Selector7~5_combout ),
	.cin(gnd),
	.combout(\Selector7~6_combout ),
	.cout());
defparam \Selector7~6 .lut_mask = 16'hFFFE;
defparam \Selector7~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector9~0 (
	.dataa(\sig_dgwb_state.s_write_mtp~q ),
	.datab(\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(gnd),
	.datad(\Selector7~6_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hEEFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_state.s_write_01_pairs (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_01_pairs~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_01_pairs .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_01_pairs .power_up = "low";

cycloneiii_lcell_comb \Selector67~2 (
	.dataa(\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datab(\Selector67~1_combout ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_01_pairs~q ),
	.cin(gnd),
	.combout(\Selector67~2_combout ),
	.cout());
defparam \Selector67~2 .lut_mask = 16'hAACC;
defparam \Selector67~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector67~3 (
	.dataa(\sig_dgwb_last_state.s_write_zeros~q ),
	.datab(\Selector67~2_combout ),
	.datac(\sig_dgwb_state.s_write_zeros~q ),
	.datad(\sig_dgwb_state.s_write_ones~q ),
	.cin(gnd),
	.combout(\Selector67~3_combout ),
	.cout());
defparam \Selector67~3 .lut_mask = 16'hACFF;
defparam \Selector67~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector67~4 (
	.dataa(\generate_wdata~q ),
	.datab(\Selector67~0_combout ),
	.datac(\Selector67~3_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector67~4_combout ),
	.cout());
defparam \Selector67~4 .lut_mask = 16'h5F3F;
defparam \Selector67~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~1 (
	.dataa(\sig_dgwb_last_state.s_write_wlat~q ),
	.datab(\sig_dgwb_state.s_write_wlat~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~1_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~1 .lut_mask = 16'hEEEE;
defparam \sig_addr_cmd[0].addr[5]~1 .sum_lutc_input = "datac";

dffeas generate_wdata(
	.clk(clk),
	.d(\sig_addr_cmd[0].addr[5]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\generate_wdata~q ),
	.prn(vcc));
defparam generate_wdata.is_wysiwyg = "true";
defparam generate_wdata.power_up = "low";

cycloneiii_lcell_comb \ac_handshake_proc~11 (
	.dataa(\sig_dgwb_state.s_idle~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_release_admin~q ),
	.cin(gnd),
	.combout(\ac_handshake_proc~11_combout ),
	.cout());
defparam \ac_handshake_proc~11 .lut_mask = 16'hAAFF;
defparam \ac_handshake_proc~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_write_block:sig_count[2]~3 (
	.dataa(\sig_addr_cmd[0].addr[5]~1_combout ),
	.datab(\generate_wdata~q ),
	.datac(\Selector12~1_combout ),
	.datad(\ac_handshake_proc~11_combout ),
	.cin(gnd),
	.combout(\ac_write_block:sig_count[2]~3_combout ),
	.cout());
defparam \ac_write_block:sig_count[2]~3 .lut_mask = 16'hFFFD;
defparam \ac_write_block:sig_count[2]~3 .sum_lutc_input = "datac";

dffeas \ac_write_block:sig_count[2] (
	.clk(clk),
	.d(\ac_write_block:sig_count[2]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[2]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[2] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[2] .power_up = "low";

dffeas \ac_write_block:sig_count[0] (
	.clk(clk),
	.d(\ac_write_block:sig_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[0]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[0] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[0] .power_up = "low";

dffeas \ac_write_block:sig_count[1] (
	.clk(clk),
	.d(\ac_write_block:sig_count[1]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[1]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[1] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[1] .power_up = "low";

cycloneiii_lcell_comb \Selector75~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ac_write_block:sig_count[0]~q ),
	.datad(\ac_write_block:sig_count[1]~q ),
	.cin(gnd),
	.combout(\Selector75~6_combout ),
	.cout());
defparam \Selector75~6 .lut_mask = 16'h0FFF;
defparam \Selector75~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_write_block:sig_count[3]~1 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[2]~2 ),
	.combout(\ac_write_block:sig_count[3]~1_combout ),
	.cout(\ac_write_block:sig_count[3]~2 ));
defparam \ac_write_block:sig_count[3]~1 .lut_mask = 16'h5A5F;
defparam \ac_write_block:sig_count[3]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \ac_write_block:sig_count[4]~1 (
	.dataa(\ac_write_block:sig_count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[3]~2 ),
	.combout(\ac_write_block:sig_count[4]~1_combout ),
	.cout(\ac_write_block:sig_count[4]~2 ));
defparam \ac_write_block:sig_count[4]~1 .lut_mask = 16'h5AAF;
defparam \ac_write_block:sig_count[4]~1 .sum_lutc_input = "cin";

dffeas \ac_write_block:sig_count[4] (
	.clk(clk),
	.d(\ac_write_block:sig_count[4]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[4]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[4] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[4] .power_up = "low";

cycloneiii_lcell_comb \ac_write_block:sig_count[5]~1 (
	.dataa(\ac_write_block:sig_count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[4]~2 ),
	.combout(\ac_write_block:sig_count[5]~1_combout ),
	.cout(\ac_write_block:sig_count[5]~2 ));
defparam \ac_write_block:sig_count[5]~1 .lut_mask = 16'h5A5F;
defparam \ac_write_block:sig_count[5]~1 .sum_lutc_input = "cin";

cycloneiii_lcell_comb \ac_write_block:sig_count[6]~1 (
	.dataa(\ac_write_block:sig_count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ac_write_block:sig_count[5]~2 ),
	.combout(\ac_write_block:sig_count[6]~1_combout ),
	.cout(\ac_write_block:sig_count[6]~2 ));
defparam \ac_write_block:sig_count[6]~1 .lut_mask = 16'h5AAF;
defparam \ac_write_block:sig_count[6]~1 .sum_lutc_input = "cin";

dffeas \ac_write_block:sig_count[6] (
	.clk(clk),
	.d(\ac_write_block:sig_count[6]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[6]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[6] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[6] .power_up = "low";

cycloneiii_lcell_comb \Equal1~0 (
	.dataa(\Selector75~5_combout ),
	.datab(\Selector75~6_combout ),
	.datac(\ac_write_block:sig_count[4]~q ),
	.datad(\ac_write_block:sig_count[6]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal0~0 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\ac_write_block:sig_count[2]~q ),
	.datac(gnd),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector26~0 (
	.dataa(\Equal1~1_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\sig_dgwb_state.s_write_zeros~q ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
defparam \Selector26~0 .lut_mask = 16'hFAFC;
defparam \Selector26~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector26~1 (
	.dataa(\sig_dgwb_state.s_write_0011_step~q ),
	.datab(\Selector26~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
defparam \Selector26~1 .lut_mask = 16'hEEEE;
defparam \Selector26~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~0 (
	.dataa(\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(\Equal0~0_combout ),
	.datac(gnd),
	.datad(\sig_dgwb_last_state.s_write_01_pairs~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~0_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~0 .lut_mask = 16'hEEFF;
defparam \sig_addr_cmd[0].addr[5]~0 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_write_zeros (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_zeros~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_zeros~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_zeros .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_zeros .power_up = "low";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~2 (
	.dataa(\sig_dgwb_last_state.s_write_0011_step~q ),
	.datab(\sig_dgwb_state.s_write_0011_step~q ),
	.datac(\sig_dgwb_state.s_write_zeros~q ),
	.datad(\sig_dgwb_last_state.s_write_zeros~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~2_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~2 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd[0].addr[5]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~3 (
	.dataa(\sig_addr_cmd[0].addr[5]~1_combout ),
	.datab(\sig_addr_cmd[0].addr[5]~2_combout ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\sig_dgwb_last_state.s_write_ones~q ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~3_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~3 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd[0].addr[5]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~4 (
	.dataa(\sig_dgwb_last_state.s_write_1100_step~q ),
	.datab(\sig_dgwb_state.s_write_1100_step~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~4_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~4 .lut_mask = 16'hEEEE;
defparam \sig_addr_cmd[0].addr[5]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~5 (
	.dataa(\sig_dgwb_state.s_release_admin~q ),
	.datab(\sig_addr_cmd[0].addr[5]~3_combout ),
	.datac(\sig_addr_cmd[0].addr[5]~4_combout ),
	.datad(\Selector12~1_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~5_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~5 .lut_mask = 16'hFEFF;
defparam \sig_addr_cmd[0].addr[5]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd~518 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\ac_write_block:sig_count[2]~q ),
	.datac(gnd),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd~518_combout ),
	.cout());
defparam \sig_addr_cmd~518 .lut_mask = 16'hEEFF;
defparam \sig_addr_cmd~518 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Equal4~0 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\ac_write_block:sig_count[2]~q ),
	.datac(\Equal1~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'hFEFE;
defparam \Equal4~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~6 (
	.dataa(\sig_dgwb_state.s_write_ones~q ),
	.datab(\sig_dgwb_state.s_write_zeros~q ),
	.datac(gnd),
	.datad(\Equal4~0_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~6_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~6 .lut_mask = 16'hEEFF;
defparam \sig_addr_cmd[0].addr[5]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \sig_addr_cmd[0].addr[5]~7 (
	.dataa(\sig_addr_cmd[0].addr[5]~0_combout ),
	.datab(\sig_addr_cmd[0].addr[5]~5_combout ),
	.datac(\sig_addr_cmd~518_combout ),
	.datad(\sig_addr_cmd[0].addr[5]~6_combout ),
	.cin(gnd),
	.combout(\sig_addr_cmd[0].addr[5]~7_combout ),
	.cout());
defparam \sig_addr_cmd[0].addr[5]~7 .lut_mask = 16'h7FFF;
defparam \sig_addr_cmd[0].addr[5]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector25~0 (
	.dataa(\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(\sig_addr_cmd~518_combout ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\sig_dgwb_state.s_write_zeros~q ),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
defparam \Selector25~0 .lut_mask = 16'hFAFC;
defparam \Selector25~0 .sum_lutc_input = "datac";

dffeas \ac_write_block:sig_count[3] (
	.clk(clk),
	.d(\ac_write_block:sig_count[3]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[3]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[3] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[3] .power_up = "low";

cycloneiii_lcell_comb \Equal1~1 (
	.dataa(\ac_write_block:sig_count[2]~q ),
	.datab(\Equal1~0_combout ),
	.datac(gnd),
	.datad(\ac_write_block:sig_count[3]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hEEFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector24~0 (
	.dataa(\Equal0~0_combout ),
	.datab(\sig_dgwb_state.s_write_zeros~q ),
	.datac(\Equal1~1_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
defparam \Selector24~0 .lut_mask = 16'hEFFF;
defparam \Selector24~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector23~0 (
	.dataa(\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(\Equal0~0_combout ),
	.datac(\sig_dgwb_state.s_write_ones~q ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
defparam \Selector23~0 .lut_mask = 16'hFEFF;
defparam \Selector23~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector58~0 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(\sig_dgwb_state.s_write_ones~q ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_0011_step~q ),
	.cin(gnd),
	.combout(\Selector58~0_combout ),
	.cout());
defparam \Selector58~0 .lut_mask = 16'hAACC;
defparam \Selector58~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgwb_wdata[24]~9 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(\Selector58~0_combout ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_1100_step~q ),
	.cin(gnd),
	.combout(\dgwb_wdata[24]~9_combout ),
	.cout());
defparam \dgwb_wdata[24]~9 .lut_mask = 16'hCC55;
defparam \dgwb_wdata[24]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgwb_wdata~11 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(\generate_wdata~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dgwb_wdata~11_combout ),
	.cout());
defparam \dgwb_wdata~11 .lut_mask = 16'hEEEE;
defparam \dgwb_wdata~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector66~0 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(\sig_dgwb_state.s_write_ones~q ),
	.datac(\sig_dgwb_state.s_write_01_pairs~q ),
	.datad(\sig_dgwb_state.s_write_0011_step~q ),
	.cin(gnd),
	.combout(\Selector66~0_combout ),
	.cout());
defparam \Selector66~0 .lut_mask = 16'hFAFC;
defparam \Selector66~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgwb_wdata[8]~10 (
	.dataa(\ac_write_block:sig_count[0]~q ),
	.datab(\Selector66~0_combout ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_1100_step~q ),
	.cin(gnd),
	.combout(\dgwb_wdata[8]~10_combout ),
	.cout());
defparam \dgwb_wdata[8]~10 .lut_mask = 16'hCC55;
defparam \dgwb_wdata[8]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \dgwb_dqs_burst~0 (
	.dataa(\sig_dgwb_state.s_wait_admin~q ),
	.datab(\sig_dgwb_state.s_release_admin~q ),
	.datac(\Selector12~0_combout ),
	.datad(\sig_dgwb_state.s_idle~q ),
	.cin(gnd),
	.combout(\dgwb_dqs_burst~0_combout ),
	.cout());
defparam \dgwb_dqs_burst~0 .lut_mask = 16'hFFF7;
defparam \dgwb_dqs_burst~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector6~0 (
	.dataa(\sig_dgwb_state.s_write_zeros~q ),
	.datab(\sig_dgwb_last_state.s_write_zeros~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hEEEE;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~0 (
	.dataa(\sig_addr_cmd~518_combout ),
	.datab(\Selector67~0_combout ),
	.datac(\Equal4~0_combout ),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(\Selector50~0_combout ),
	.cout());
defparam \Selector50~0 .lut_mask = 16'hBFFF;
defparam \Selector50~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~2 (
	.dataa(\Selector50~1_combout ),
	.datab(\sig_dgwb_last_state.s_write_wlat~q ),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector50~2_combout ),
	.cout());
defparam \Selector50~2 .lut_mask = 16'hEEFF;
defparam \Selector50~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector50~3 (
	.dataa(\Selector50~0_combout ),
	.datab(\Selector50~2_combout ),
	.datac(\Equal0~0_combout ),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\Selector50~3_combout ),
	.cout());
defparam \Selector50~3 .lut_mask = 16'hFF7F;
defparam \Selector50~3 .sum_lutc_input = "datac";

dffeas \sig_dgwb_last_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgwb_state.s_release_admin~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_release_admin .power_up = "low";

cycloneiii_lcell_comb \ac_handshake_proc~2 (
	.dataa(\sig_dgwb_last_state.s_release_admin~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sig_dgwb_state.s_idle~q ),
	.cin(gnd),
	.combout(\ac_handshake_proc~2_combout ),
	.cout());
defparam \ac_handshake_proc~2 .lut_mask = 16'hAAFF;
defparam \ac_handshake_proc~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector57~0 (
	.dataa(\ac_write_block:sig_count[1]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector57~0_combout ),
	.cout());
defparam \Selector57~0 .lut_mask = 16'hFAFC;
defparam \Selector57~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector65~0 (
	.dataa(\ac_write_block:sig_count[1]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector65~0_combout ),
	.cout());
defparam \Selector65~0 .lut_mask = 16'hFAFC;
defparam \Selector65~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector56~0 (
	.dataa(\ac_write_block:sig_count[2]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector56~0_combout ),
	.cout());
defparam \Selector56~0 .lut_mask = 16'hFAFC;
defparam \Selector56~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector64~0 (
	.dataa(\ac_write_block:sig_count[2]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector64~0_combout ),
	.cout());
defparam \Selector64~0 .lut_mask = 16'hFAFC;
defparam \Selector64~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector55~0 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector55~0_combout ),
	.cout());
defparam \Selector55~0 .lut_mask = 16'hFAFC;
defparam \Selector55~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector63~0 (
	.dataa(\ac_write_block:sig_count[3]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector63~0_combout ),
	.cout());
defparam \Selector63~0 .lut_mask = 16'hFAFC;
defparam \Selector63~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector54~3 (
	.dataa(\ac_write_block:sig_count[4]~q ),
	.datab(\sig_dgwb_state.s_write_wlat~q ),
	.datac(\generate_wdata~q ),
	.datad(\dgwb_wdata[24]~9_combout ),
	.cin(gnd),
	.combout(\Selector54~3_combout ),
	.cout());
defparam \Selector54~3 .lut_mask = 16'hFFB8;
defparam \Selector54~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector62~2 (
	.dataa(\ac_write_block:sig_count[4]~q ),
	.datab(\sig_dgwb_state.s_write_wlat~q ),
	.datac(\generate_wdata~q ),
	.datad(\dgwb_wdata[8]~10_combout ),
	.cin(gnd),
	.combout(\Selector62~2_combout ),
	.cout());
defparam \Selector62~2 .lut_mask = 16'hFFB8;
defparam \Selector62~2 .sum_lutc_input = "datac";

dffeas \ac_write_block:sig_count[5] (
	.clk(clk),
	.d(\ac_write_block:sig_count[5]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[5]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[5] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[5] .power_up = "low";

cycloneiii_lcell_comb \Selector53~0 (
	.dataa(\ac_write_block:sig_count[5]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector53~0_combout ),
	.cout());
defparam \Selector53~0 .lut_mask = 16'hFAFC;
defparam \Selector53~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector61~0 (
	.dataa(\ac_write_block:sig_count[5]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector61~0_combout ),
	.cout());
defparam \Selector61~0 .lut_mask = 16'hFAFC;
defparam \Selector61~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector52~0 (
	.dataa(\ac_write_block:sig_count[6]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector52~0_combout ),
	.cout());
defparam \Selector52~0 .lut_mask = 16'hFAFC;
defparam \Selector52~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector60~0 (
	.dataa(\ac_write_block:sig_count[6]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector60~0_combout ),
	.cout());
defparam \Selector60~0 .lut_mask = 16'hFAFC;
defparam \Selector60~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \ac_write_block:sig_count[7]~1 (
	.dataa(\ac_write_block:sig_count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ac_write_block:sig_count[6]~2 ),
	.combout(\ac_write_block:sig_count[7]~1_combout ),
	.cout());
defparam \ac_write_block:sig_count[7]~1 .lut_mask = 16'h5A5A;
defparam \ac_write_block:sig_count[7]~1 .sum_lutc_input = "cin";

dffeas \ac_write_block:sig_count[7] (
	.clk(clk),
	.d(\ac_write_block:sig_count[7]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\Selector67~4_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[2]~3_combout ),
	.q(\ac_write_block:sig_count[7]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[7] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[7] .power_up = "low";

cycloneiii_lcell_comb \Selector51~0 (
	.dataa(\ac_write_block:sig_count[7]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[24]~9_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector51~0_combout ),
	.cout());
defparam \Selector51~0 .lut_mask = 16'hFAFC;
defparam \Selector51~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \Selector59~0 (
	.dataa(\ac_write_block:sig_count[7]~q ),
	.datab(\generate_wdata~q ),
	.datac(\dgwb_wdata[8]~10_combout ),
	.datad(\sig_dgwb_state.s_write_wlat~q ),
	.cin(gnd),
	.combout(\Selector59~0_combout ),
	.cout());
defparam \Selector59~0 .lut_mask = 16'hFAFC;
defparam \Selector59~0 .sum_lutc_input = "datac";

endmodule

module altera_ddr_altera_ddr_phy_alt_mem_phy_write_dp_fr (
	phy_clk_1x,
	q_b_34,
	q_b_32,
	q_b_35,
	q_b_33,
	q_b_16,
	dgwb_wdata_24,
	q_b_0,
	dgwb_wdata_8,
	q_b_17,
	q_b_1,
	q_b_18,
	q_b_2,
	q_b_19,
	q_b_3,
	q_b_20,
	q_b_4,
	q_b_21,
	q_b_5,
	q_b_22,
	q_b_6,
	q_b_23,
	q_b_7,
	q_b_24,
	q_b_8,
	q_b_25,
	q_b_9,
	q_b_26,
	q_b_10,
	q_b_27,
	q_b_11,
	q_b_28,
	q_b_12,
	q_b_29,
	q_b_13,
	q_b_30,
	q_b_14,
	q_b_31,
	q_b_15,
	reset_phy_clk_1x_n,
	ctl_init_success,
	wdp_dm_l_2x_0,
	wdp_dm_h_2x_0,
	wdp_dm_l_2x_1,
	wdp_dm_h_2x_1,
	control_wlat_r_0,
	control_doing_wr,
	Equal6,
	control_doing_wr1,
	control_doing_wr2,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	wdp_wdata_l_2x_0,
	wdp_wdata_h_2x_0,
	dq_oe_2x_0,
	wdp_wdata_l_2x_1,
	wdp_wdata_h_2x_1,
	wdp_wdata_l_2x_2,
	wdp_wdata_h_2x_2,
	wdp_wdata_l_2x_3,
	wdp_wdata_h_2x_3,
	wdp_wdata_l_2x_4,
	wdp_wdata_h_2x_4,
	dq_oe_2x_1,
	wdp_wdata_l_2x_5,
	wdp_wdata_h_2x_5,
	wdp_wdata_l_2x_6,
	wdp_wdata_h_2x_6,
	wdp_wdata_l_2x_7,
	wdp_wdata_h_2x_7,
	wdp_wdata_l_2x_8,
	wdp_wdata_h_2x_8,
	dq_oe_2x_2,
	wdp_wdata_l_2x_9,
	wdp_wdata_h_2x_9,
	wdp_wdata_l_2x_10,
	wdp_wdata_h_2x_10,
	wdp_wdata_l_2x_11,
	wdp_wdata_h_2x_11,
	wdp_wdata_l_2x_12,
	wdp_wdata_h_2x_12,
	dq_oe_2x_3,
	wdp_wdata_l_2x_13,
	wdp_wdata_h_2x_13,
	wdp_wdata_l_2x_14,
	wdp_wdata_h_2x_14,
	wdp_wdata_l_2x_15,
	wdp_wdata_h_2x_15,
	wdp_wdqs_2x_1,
	wdp_wdqs_oe_2x_0,
	dgwb_wdata_25,
	dgwb_wdata_9,
	dgwb_wdata_26,
	dgwb_wdata_10,
	dgwb_wdata_27,
	dgwb_wdata_11,
	dgwb_wdata_28,
	dgwb_wdata_12,
	dgwb_wdata_29,
	dgwb_wdata_13,
	dgwb_wdata_30,
	dgwb_wdata_14,
	dgwb_wdata_31,
	dgwb_wdata_15,
	control_dqs_burst_0,
	dqs_burst_cas4,
	dqs_burst_cas3)/* synthesis synthesis_greybox=1 */;
input 	phy_clk_1x;
input 	q_b_34;
input 	q_b_32;
input 	q_b_35;
input 	q_b_33;
input 	q_b_16;
input 	dgwb_wdata_24;
input 	q_b_0;
input 	dgwb_wdata_8;
input 	q_b_17;
input 	q_b_1;
input 	q_b_18;
input 	q_b_2;
input 	q_b_19;
input 	q_b_3;
input 	q_b_20;
input 	q_b_4;
input 	q_b_21;
input 	q_b_5;
input 	q_b_22;
input 	q_b_6;
input 	q_b_23;
input 	q_b_7;
input 	q_b_24;
input 	q_b_8;
input 	q_b_25;
input 	q_b_9;
input 	q_b_26;
input 	q_b_10;
input 	q_b_27;
input 	q_b_11;
input 	q_b_28;
input 	q_b_12;
input 	q_b_29;
input 	q_b_13;
input 	q_b_30;
input 	q_b_14;
input 	q_b_31;
input 	q_b_15;
input 	reset_phy_clk_1x_n;
input 	ctl_init_success;
output 	wdp_dm_l_2x_0;
output 	wdp_dm_h_2x_0;
output 	wdp_dm_l_2x_1;
output 	wdp_dm_h_2x_1;
input 	control_wlat_r_0;
input 	control_doing_wr;
input 	Equal6;
input 	control_doing_wr1;
input 	control_doing_wr2;
input 	dgwb_wdp_ovride;
input 	seq_wdp_ovride;
output 	wdp_wdata_l_2x_0;
output 	wdp_wdata_h_2x_0;
output 	dq_oe_2x_0;
output 	wdp_wdata_l_2x_1;
output 	wdp_wdata_h_2x_1;
output 	wdp_wdata_l_2x_2;
output 	wdp_wdata_h_2x_2;
output 	wdp_wdata_l_2x_3;
output 	wdp_wdata_h_2x_3;
output 	wdp_wdata_l_2x_4;
output 	wdp_wdata_h_2x_4;
output 	dq_oe_2x_1;
output 	wdp_wdata_l_2x_5;
output 	wdp_wdata_h_2x_5;
output 	wdp_wdata_l_2x_6;
output 	wdp_wdata_h_2x_6;
output 	wdp_wdata_l_2x_7;
output 	wdp_wdata_h_2x_7;
output 	wdp_wdata_l_2x_8;
output 	wdp_wdata_h_2x_8;
output 	dq_oe_2x_2;
output 	wdp_wdata_l_2x_9;
output 	wdp_wdata_h_2x_9;
output 	wdp_wdata_l_2x_10;
output 	wdp_wdata_h_2x_10;
output 	wdp_wdata_l_2x_11;
output 	wdp_wdata_h_2x_11;
output 	wdp_wdata_l_2x_12;
output 	wdp_wdata_h_2x_12;
output 	dq_oe_2x_3;
output 	wdp_wdata_l_2x_13;
output 	wdp_wdata_h_2x_13;
output 	wdp_wdata_l_2x_14;
output 	wdp_wdata_h_2x_14;
output 	wdp_wdata_l_2x_15;
output 	wdp_wdata_h_2x_15;
output 	wdp_wdqs_2x_1;
output 	wdp_wdqs_oe_2x_0;
input 	dgwb_wdata_25;
input 	dgwb_wdata_9;
input 	dgwb_wdata_26;
input 	dgwb_wdata_10;
input 	dgwb_wdata_27;
input 	dgwb_wdata_11;
input 	dgwb_wdata_28;
input 	dgwb_wdata_12;
input 	dgwb_wdata_29;
input 	dgwb_wdata_13;
input 	dgwb_wdata_30;
input 	dgwb_wdata_14;
input 	dgwb_wdata_31;
input 	dgwb_wdata_15;
input 	control_dqs_burst_0;
input 	dqs_burst_cas4;
input 	dqs_burst_cas3;

wire gnd;
wire vcc;

assign gnd = 1'b0;
assign vcc = 1'b1;

wire \wdp_dm_l_2x~2_combout ;
wire \wdp_dm_h_2x~2_combout ;
wire \wdp_dm_l_2x~3_combout ;
wire \wdp_dm_h_2x~3_combout ;
wire \mem_wdata[16]~0_combout ;
wire \mem_wdata[0]~1_combout ;
wire \mem_wdata_valid[0]~0_combout ;
wire \mem_wdata[17]~2_combout ;
wire \mem_wdata[1]~3_combout ;
wire \mem_wdata[18]~4_combout ;
wire \mem_wdata[2]~5_combout ;
wire \mem_wdata[19]~6_combout ;
wire \mem_wdata[3]~7_combout ;
wire \mem_wdata[20]~8_combout ;
wire \mem_wdata[4]~9_combout ;
wire \mem_wdata[21]~10_combout ;
wire \mem_wdata[5]~11_combout ;
wire \mem_wdata[22]~12_combout ;
wire \mem_wdata[6]~13_combout ;
wire \mem_wdata[23]~14_combout ;
wire \mem_wdata[7]~15_combout ;
wire \mem_wdata[24]~16_combout ;
wire \mem_wdata[8]~17_combout ;
wire \mem_wdata[25]~18_combout ;
wire \mem_wdata[9]~19_combout ;
wire \mem_wdata[26]~20_combout ;
wire \mem_wdata[10]~21_combout ;
wire \mem_wdata[27]~22_combout ;
wire \mem_wdata[11]~23_combout ;
wire \mem_wdata[28]~24_combout ;
wire \mem_wdata[12]~25_combout ;
wire \mem_wdata[29]~26_combout ;
wire \mem_wdata[13]~27_combout ;
wire \mem_wdata[30]~28_combout ;
wire \mem_wdata[14]~29_combout ;
wire \mem_wdata[31]~30_combout ;
wire \mem_wdata[15]~31_combout ;
wire \mem_dqs_burst[0]~0_combout ;
wire \mem_dqs_burst[0]~1_combout ;


dffeas \wdp_dm_l_2x[0] (
	.clk(phy_clk_1x),
	.d(\wdp_dm_l_2x~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_dm_l_2x_0),
	.prn(vcc));
defparam \wdp_dm_l_2x[0] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[0] .power_up = "low";

dffeas \wdp_dm_h_2x[0] (
	.clk(phy_clk_1x),
	.d(\wdp_dm_h_2x~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_dm_h_2x_0),
	.prn(vcc));
defparam \wdp_dm_h_2x[0] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[0] .power_up = "low";

dffeas \wdp_dm_l_2x[1] (
	.clk(phy_clk_1x),
	.d(\wdp_dm_l_2x~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_dm_l_2x_1),
	.prn(vcc));
defparam \wdp_dm_l_2x[1] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[1] .power_up = "low";

dffeas \wdp_dm_h_2x[1] (
	.clk(phy_clk_1x),
	.d(\wdp_dm_h_2x~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_dm_h_2x_1),
	.prn(vcc));
defparam \wdp_dm_h_2x[1] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[1] .power_up = "low";

dffeas \wdp_wdata_l_2x[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[16]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_0),
	.prn(vcc));
defparam \wdp_wdata_l_2x[0] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[0] .power_up = "low";

dffeas \wdp_wdata_h_2x[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_0),
	.prn(vcc));
defparam \wdp_wdata_h_2x[0] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[0] .power_up = "low";

dffeas \dq_oe_2x[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dq_oe_2x_0),
	.prn(vcc));
defparam \dq_oe_2x[0] .is_wysiwyg = "true";
defparam \dq_oe_2x[0] .power_up = "low";

dffeas \wdp_wdata_l_2x[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[17]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_1),
	.prn(vcc));
defparam \wdp_wdata_l_2x[1] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[1] .power_up = "low";

dffeas \wdp_wdata_h_2x[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_1),
	.prn(vcc));
defparam \wdp_wdata_h_2x[1] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[1] .power_up = "low";

dffeas \wdp_wdata_l_2x[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[18]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_2),
	.prn(vcc));
defparam \wdp_wdata_l_2x[2] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[2] .power_up = "low";

dffeas \wdp_wdata_h_2x[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[2]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_2),
	.prn(vcc));
defparam \wdp_wdata_h_2x[2] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[2] .power_up = "low";

dffeas \wdp_wdata_l_2x[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[19]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_3),
	.prn(vcc));
defparam \wdp_wdata_l_2x[3] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[3] .power_up = "low";

dffeas \wdp_wdata_h_2x[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[3]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_3),
	.prn(vcc));
defparam \wdp_wdata_h_2x[3] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[3] .power_up = "low";

dffeas \wdp_wdata_l_2x[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[20]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_4),
	.prn(vcc));
defparam \wdp_wdata_l_2x[4] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[4] .power_up = "low";

dffeas \wdp_wdata_h_2x[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[4]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_4),
	.prn(vcc));
defparam \wdp_wdata_h_2x[4] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[4] .power_up = "low";

dffeas \dq_oe_2x[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dq_oe_2x_1),
	.prn(vcc));
defparam \dq_oe_2x[1] .is_wysiwyg = "true";
defparam \dq_oe_2x[1] .power_up = "low";

dffeas \wdp_wdata_l_2x[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[21]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_5),
	.prn(vcc));
defparam \wdp_wdata_l_2x[5] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[5] .power_up = "low";

dffeas \wdp_wdata_h_2x[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[5]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_5),
	.prn(vcc));
defparam \wdp_wdata_h_2x[5] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[5] .power_up = "low";

dffeas \wdp_wdata_l_2x[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[22]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_6),
	.prn(vcc));
defparam \wdp_wdata_l_2x[6] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[6] .power_up = "low";

dffeas \wdp_wdata_h_2x[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[6]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_6),
	.prn(vcc));
defparam \wdp_wdata_h_2x[6] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[6] .power_up = "low";

dffeas \wdp_wdata_l_2x[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[23]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_7),
	.prn(vcc));
defparam \wdp_wdata_l_2x[7] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[7] .power_up = "low";

dffeas \wdp_wdata_h_2x[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[7]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_7),
	.prn(vcc));
defparam \wdp_wdata_h_2x[7] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[7] .power_up = "low";

dffeas \wdp_wdata_l_2x[8] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[24]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_8),
	.prn(vcc));
defparam \wdp_wdata_l_2x[8] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[8] .power_up = "low";

dffeas \wdp_wdata_h_2x[8] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[8]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_8),
	.prn(vcc));
defparam \wdp_wdata_h_2x[8] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[8] .power_up = "low";

dffeas \dq_oe_2x[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dq_oe_2x_2),
	.prn(vcc));
defparam \dq_oe_2x[2] .is_wysiwyg = "true";
defparam \dq_oe_2x[2] .power_up = "low";

dffeas \wdp_wdata_l_2x[9] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[25]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_9),
	.prn(vcc));
defparam \wdp_wdata_l_2x[9] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[9] .power_up = "low";

dffeas \wdp_wdata_h_2x[9] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[9]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_9),
	.prn(vcc));
defparam \wdp_wdata_h_2x[9] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[9] .power_up = "low";

dffeas \wdp_wdata_l_2x[10] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[26]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_10),
	.prn(vcc));
defparam \wdp_wdata_l_2x[10] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[10] .power_up = "low";

dffeas \wdp_wdata_h_2x[10] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[10]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_10),
	.prn(vcc));
defparam \wdp_wdata_h_2x[10] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[10] .power_up = "low";

dffeas \wdp_wdata_l_2x[11] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[27]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_11),
	.prn(vcc));
defparam \wdp_wdata_l_2x[11] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[11] .power_up = "low";

dffeas \wdp_wdata_h_2x[11] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[11]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_11),
	.prn(vcc));
defparam \wdp_wdata_h_2x[11] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[11] .power_up = "low";

dffeas \wdp_wdata_l_2x[12] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[28]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_12),
	.prn(vcc));
defparam \wdp_wdata_l_2x[12] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[12] .power_up = "low";

dffeas \wdp_wdata_h_2x[12] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[12]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_12),
	.prn(vcc));
defparam \wdp_wdata_h_2x[12] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[12] .power_up = "low";

dffeas \dq_oe_2x[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dq_oe_2x_3),
	.prn(vcc));
defparam \dq_oe_2x[3] .is_wysiwyg = "true";
defparam \dq_oe_2x[3] .power_up = "low";

dffeas \wdp_wdata_l_2x[13] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[29]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_13),
	.prn(vcc));
defparam \wdp_wdata_l_2x[13] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[13] .power_up = "low";

dffeas \wdp_wdata_h_2x[13] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[13]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_13),
	.prn(vcc));
defparam \wdp_wdata_h_2x[13] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[13] .power_up = "low";

dffeas \wdp_wdata_l_2x[14] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[30]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_14),
	.prn(vcc));
defparam \wdp_wdata_l_2x[14] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[14] .power_up = "low";

dffeas \wdp_wdata_h_2x[14] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[14]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_14),
	.prn(vcc));
defparam \wdp_wdata_h_2x[14] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[14] .power_up = "low";

dffeas \wdp_wdata_l_2x[15] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[31]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_l_2x_15),
	.prn(vcc));
defparam \wdp_wdata_l_2x[15] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[15] .power_up = "low";

dffeas \wdp_wdata_h_2x[15] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[15]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdata_h_2x_15),
	.prn(vcc));
defparam \wdp_wdata_h_2x[15] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[15] .power_up = "low";

dffeas \wdp_wdqs_2x[1] (
	.clk(phy_clk_1x),
	.d(wdp_wdqs_oe_2x_0),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdqs_2x_1),
	.prn(vcc));
defparam \wdp_wdqs_2x[1] .is_wysiwyg = "true";
defparam \wdp_wdqs_2x[1] .power_up = "low";

dffeas \wdp_wdqs_oe_2x[0] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wdp_wdqs_oe_2x_0),
	.prn(vcc));
defparam \wdp_wdqs_oe_2x[0] .is_wysiwyg = "true";
defparam \wdp_wdqs_oe_2x[0] .power_up = "low";

cycloneiii_lcell_comb \wdp_dm_l_2x~2 (
	.dataa(control_doing_wr1),
	.datab(control_doing_wr2),
	.datac(q_b_34),
	.datad(seq_wdp_ovride),
	.cin(gnd),
	.combout(\wdp_dm_l_2x~2_combout ),
	.cout());
defparam \wdp_dm_l_2x~2 .lut_mask = 16'h7FFF;
defparam \wdp_dm_l_2x~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdp_dm_h_2x~2 (
	.dataa(control_doing_wr1),
	.datab(control_doing_wr2),
	.datac(q_b_32),
	.datad(seq_wdp_ovride),
	.cin(gnd),
	.combout(\wdp_dm_h_2x~2_combout ),
	.cout());
defparam \wdp_dm_h_2x~2 .lut_mask = 16'h7FFF;
defparam \wdp_dm_h_2x~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdp_dm_l_2x~3 (
	.dataa(control_doing_wr1),
	.datab(control_doing_wr2),
	.datac(q_b_35),
	.datad(seq_wdp_ovride),
	.cin(gnd),
	.combout(\wdp_dm_l_2x~3_combout ),
	.cout());
defparam \wdp_dm_l_2x~3 .lut_mask = 16'h7FFF;
defparam \wdp_dm_l_2x~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \wdp_dm_h_2x~3 (
	.dataa(control_doing_wr1),
	.datab(control_doing_wr2),
	.datac(q_b_33),
	.datad(seq_wdp_ovride),
	.cin(gnd),
	.combout(\wdp_dm_h_2x~3_combout ),
	.cout());
defparam \wdp_dm_h_2x~3 .lut_mask = 16'h7FFF;
defparam \wdp_dm_h_2x~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[16]~0 (
	.dataa(q_b_16),
	.datab(dgwb_wdata_24),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[16]~0_combout ),
	.cout());
defparam \mem_wdata[16]~0 .lut_mask = 16'hEFFE;
defparam \mem_wdata[16]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[0]~1 (
	.dataa(q_b_0),
	.datab(dgwb_wdata_8),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[0]~1_combout ),
	.cout());
defparam \mem_wdata[0]~1 .lut_mask = 16'hEFFE;
defparam \mem_wdata[0]~1 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata_valid[0]~0 (
	.dataa(control_doing_wr1),
	.datab(control_doing_wr2),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata_valid[0]~0_combout ),
	.cout());
defparam \mem_wdata_valid[0]~0 .lut_mask = 16'hFEFF;
defparam \mem_wdata_valid[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[17]~2 (
	.dataa(q_b_17),
	.datab(dgwb_wdata_25),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[17]~2_combout ),
	.cout());
defparam \mem_wdata[17]~2 .lut_mask = 16'hEFFE;
defparam \mem_wdata[17]~2 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[1]~3 (
	.dataa(q_b_1),
	.datab(dgwb_wdata_9),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[1]~3_combout ),
	.cout());
defparam \mem_wdata[1]~3 .lut_mask = 16'hEFFE;
defparam \mem_wdata[1]~3 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[18]~4 (
	.dataa(q_b_18),
	.datab(dgwb_wdata_26),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[18]~4_combout ),
	.cout());
defparam \mem_wdata[18]~4 .lut_mask = 16'hEFFE;
defparam \mem_wdata[18]~4 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[2]~5 (
	.dataa(q_b_2),
	.datab(dgwb_wdata_10),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[2]~5_combout ),
	.cout());
defparam \mem_wdata[2]~5 .lut_mask = 16'hEFFE;
defparam \mem_wdata[2]~5 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[19]~6 (
	.dataa(q_b_19),
	.datab(dgwb_wdata_27),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[19]~6_combout ),
	.cout());
defparam \mem_wdata[19]~6 .lut_mask = 16'hEFFE;
defparam \mem_wdata[19]~6 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[3]~7 (
	.dataa(q_b_3),
	.datab(dgwb_wdata_11),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[3]~7_combout ),
	.cout());
defparam \mem_wdata[3]~7 .lut_mask = 16'hEFFE;
defparam \mem_wdata[3]~7 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[20]~8 (
	.dataa(q_b_20),
	.datab(dgwb_wdata_28),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[20]~8_combout ),
	.cout());
defparam \mem_wdata[20]~8 .lut_mask = 16'hEFFE;
defparam \mem_wdata[20]~8 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[4]~9 (
	.dataa(q_b_4),
	.datab(dgwb_wdata_12),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[4]~9_combout ),
	.cout());
defparam \mem_wdata[4]~9 .lut_mask = 16'hEFFE;
defparam \mem_wdata[4]~9 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[21]~10 (
	.dataa(q_b_21),
	.datab(dgwb_wdata_29),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[21]~10_combout ),
	.cout());
defparam \mem_wdata[21]~10 .lut_mask = 16'hEFFE;
defparam \mem_wdata[21]~10 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[5]~11 (
	.dataa(q_b_5),
	.datab(dgwb_wdata_13),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[5]~11_combout ),
	.cout());
defparam \mem_wdata[5]~11 .lut_mask = 16'hEFFE;
defparam \mem_wdata[5]~11 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[22]~12 (
	.dataa(q_b_22),
	.datab(dgwb_wdata_30),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[22]~12_combout ),
	.cout());
defparam \mem_wdata[22]~12 .lut_mask = 16'hEFFE;
defparam \mem_wdata[22]~12 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[6]~13 (
	.dataa(q_b_6),
	.datab(dgwb_wdata_14),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[6]~13_combout ),
	.cout());
defparam \mem_wdata[6]~13 .lut_mask = 16'hEFFE;
defparam \mem_wdata[6]~13 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[23]~14 (
	.dataa(q_b_23),
	.datab(dgwb_wdata_31),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[23]~14_combout ),
	.cout());
defparam \mem_wdata[23]~14 .lut_mask = 16'hEFFE;
defparam \mem_wdata[23]~14 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[7]~15 (
	.dataa(q_b_7),
	.datab(dgwb_wdata_15),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[7]~15_combout ),
	.cout());
defparam \mem_wdata[7]~15 .lut_mask = 16'hEFFE;
defparam \mem_wdata[7]~15 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[24]~16 (
	.dataa(q_b_24),
	.datab(dgwb_wdata_24),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[24]~16_combout ),
	.cout());
defparam \mem_wdata[24]~16 .lut_mask = 16'hEFFE;
defparam \mem_wdata[24]~16 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[8]~17 (
	.dataa(q_b_8),
	.datab(dgwb_wdata_8),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[8]~17_combout ),
	.cout());
defparam \mem_wdata[8]~17 .lut_mask = 16'hEFFE;
defparam \mem_wdata[8]~17 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[25]~18 (
	.dataa(q_b_25),
	.datab(dgwb_wdata_25),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[25]~18_combout ),
	.cout());
defparam \mem_wdata[25]~18 .lut_mask = 16'hEFFE;
defparam \mem_wdata[25]~18 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[9]~19 (
	.dataa(q_b_9),
	.datab(dgwb_wdata_9),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[9]~19_combout ),
	.cout());
defparam \mem_wdata[9]~19 .lut_mask = 16'hEFFE;
defparam \mem_wdata[9]~19 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[26]~20 (
	.dataa(q_b_26),
	.datab(dgwb_wdata_26),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[26]~20_combout ),
	.cout());
defparam \mem_wdata[26]~20 .lut_mask = 16'hEFFE;
defparam \mem_wdata[26]~20 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[10]~21 (
	.dataa(q_b_10),
	.datab(dgwb_wdata_10),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[10]~21_combout ),
	.cout());
defparam \mem_wdata[10]~21 .lut_mask = 16'hEFFE;
defparam \mem_wdata[10]~21 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[27]~22 (
	.dataa(q_b_27),
	.datab(dgwb_wdata_27),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[27]~22_combout ),
	.cout());
defparam \mem_wdata[27]~22 .lut_mask = 16'hEFFE;
defparam \mem_wdata[27]~22 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[11]~23 (
	.dataa(q_b_11),
	.datab(dgwb_wdata_11),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[11]~23_combout ),
	.cout());
defparam \mem_wdata[11]~23 .lut_mask = 16'hEFFE;
defparam \mem_wdata[11]~23 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[28]~24 (
	.dataa(q_b_28),
	.datab(dgwb_wdata_28),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[28]~24_combout ),
	.cout());
defparam \mem_wdata[28]~24 .lut_mask = 16'hEFFE;
defparam \mem_wdata[28]~24 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[12]~25 (
	.dataa(q_b_12),
	.datab(dgwb_wdata_12),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[12]~25_combout ),
	.cout());
defparam \mem_wdata[12]~25 .lut_mask = 16'hEFFE;
defparam \mem_wdata[12]~25 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[29]~26 (
	.dataa(q_b_29),
	.datab(dgwb_wdata_29),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[29]~26_combout ),
	.cout());
defparam \mem_wdata[29]~26 .lut_mask = 16'hEFFE;
defparam \mem_wdata[29]~26 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[13]~27 (
	.dataa(q_b_13),
	.datab(dgwb_wdata_13),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[13]~27_combout ),
	.cout());
defparam \mem_wdata[13]~27 .lut_mask = 16'hEFFE;
defparam \mem_wdata[13]~27 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[30]~28 (
	.dataa(q_b_30),
	.datab(dgwb_wdata_30),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[30]~28_combout ),
	.cout());
defparam \mem_wdata[30]~28 .lut_mask = 16'hEFFE;
defparam \mem_wdata[30]~28 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[14]~29 (
	.dataa(q_b_14),
	.datab(dgwb_wdata_14),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[14]~29_combout ),
	.cout());
defparam \mem_wdata[14]~29 .lut_mask = 16'hEFFE;
defparam \mem_wdata[14]~29 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[31]~30 (
	.dataa(q_b_31),
	.datab(dgwb_wdata_31),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[31]~30_combout ),
	.cout());
defparam \mem_wdata[31]~30 .lut_mask = 16'hEFFE;
defparam \mem_wdata[31]~30 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_wdata[15]~31 (
	.dataa(q_b_15),
	.datab(dgwb_wdata_15),
	.datac(dgwb_wdp_ovride),
	.datad(ctl_init_success),
	.cin(gnd),
	.combout(\mem_wdata[15]~31_combout ),
	.cout());
defparam \mem_wdata[15]~31 .lut_mask = 16'hEFFE;
defparam \mem_wdata[15]~31 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_dqs_burst[0]~0 (
	.dataa(dqs_burst_cas4),
	.datab(dqs_burst_cas3),
	.datac(control_wlat_r_0),
	.datad(control_doing_wr),
	.cin(gnd),
	.combout(\mem_dqs_burst[0]~0_combout ),
	.cout());
defparam \mem_dqs_burst[0]~0 .lut_mask = 16'hEFFE;
defparam \mem_dqs_burst[0]~0 .sum_lutc_input = "datac";

cycloneiii_lcell_comb \mem_dqs_burst[0]~1 (
	.dataa(seq_wdp_ovride),
	.datab(control_dqs_burst_0),
	.datac(\mem_dqs_burst[0]~0_combout ),
	.datad(Equal6),
	.cin(gnd),
	.combout(\mem_dqs_burst[0]~1_combout ),
	.cout());
defparam \mem_dqs_burst[0]~1 .lut_mask = 16'hFAFC;
defparam \mem_dqs_burst[0]~1 .sum_lutc_input = "datac";

endmodule
